VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO sram_0rw1r1w_16_256_lapis20
   CLASS BLOCK ;
   SIZE 899.4 BY 976.68 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER MET4 ;
         RECT  144.44 0.0 145.0 1.48 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER MET4 ;
         RECT  161.0 0.0 161.56 1.48 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER MET4 ;
         RECT  178.48 0.0 179.04 1.48 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER MET4 ;
         RECT  195.04 0.0 195.6 1.48 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER MET4 ;
         RECT  210.68 0.0 211.24 1.48 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER MET4 ;
         RECT  227.24 0.0 227.8 1.48 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER MET4 ;
         RECT  244.72 0.0 245.28 1.48 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER MET4 ;
         RECT  261.28 0.0 261.84 1.48 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER MET4 ;
         RECT  276.92 0.0 277.48 1.48 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER MET4 ;
         RECT  293.48 0.0 294.04 1.48 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER MET4 ;
         RECT  310.96 0.0 311.52 1.48 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER MET4 ;
         RECT  327.52 0.0 328.08 1.48 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER MET4 ;
         RECT  343.16 0.0 343.72 1.48 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER MET4 ;
         RECT  359.72 0.0 360.28 1.48 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER MET4 ;
         RECT  377.2 0.0 377.76 1.48 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER MET4 ;
         RECT  393.76 0.0 394.32 1.48 ;
      END
   END din0[15]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER MET4 ;
         RECT  112.24 0.0 112.8 1.48 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER MET4 ;
         RECT  128.8 0.0 129.36 1.48 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER MET3 ;
         RECT  0.0 295.32 1.48 295.88 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER MET3 ;
         RECT  0.0 303.6 1.48 304.16 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER MET3 ;
         RECT  0.0 310.96 1.48 311.52 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER MET3 ;
         RECT  0.0 321.08 1.48 321.64 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER MET3 ;
         RECT  0.0 328.44 1.48 329.0 ;
      END
   END addr0[6]
   PIN addr0[7]
      DIRECTION INPUT ;
      PORT
         LAYER MET3 ;
         RECT  0.0 336.72 1.48 337.28 ;
      END
   END addr0[7]
   PIN addr1[0]
      DIRECTION INPUT ;
      PORT
         LAYER MET4 ;
         RECT  770.04 975.2 770.6 976.68 ;
      END
   END addr1[0]
   PIN addr1[1]
      DIRECTION INPUT ;
      PORT
         LAYER MET4 ;
         RECT  754.4 975.2 754.96 976.68 ;
      END
   END addr1[1]
   PIN addr1[2]
      DIRECTION INPUT ;
      PORT
         LAYER MET3 ;
         RECT  897.92 88.32 899.4 88.88 ;
      END
   END addr1[2]
   PIN addr1[3]
      DIRECTION INPUT ;
      PORT
         LAYER MET3 ;
         RECT  897.92 80.04 899.4 80.6 ;
      END
   END addr1[3]
   PIN addr1[4]
      DIRECTION INPUT ;
      PORT
         LAYER MET4 ;
         RECT  821.56 0.0 822.12 1.48 ;
      END
   END addr1[4]
   PIN addr1[5]
      DIRECTION INPUT ;
      PORT
         LAYER MET4 ;
         RECT  818.8 0.0 819.36 1.48 ;
      END
   END addr1[5]
   PIN addr1[6]
      DIRECTION INPUT ;
      PORT
         LAYER MET4 ;
         RECT  820.64 0.0 821.2 1.48 ;
      END
   END addr1[6]
   PIN addr1[7]
      DIRECTION INPUT ;
      PORT
         LAYER MET4 ;
         RECT  819.72 0.0 820.28 1.48 ;
      END
   END addr1[7]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER MET3 ;
         RECT  0.0 11.96 1.48 12.52 ;
      END
   END csb0
   PIN csb1
      DIRECTION INPUT ;
      PORT
         LAYER MET3 ;
         RECT  897.92 960.48 899.4 961.04 ;
      END
   END csb1
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER MET4 ;
         RECT  36.8 0.0 37.36 1.48 ;
      END
   END clk0
   PIN clk1
      DIRECTION INPUT ;
      PORT
         LAYER MET4 ;
         RECT  862.04 975.2 862.6 976.68 ;
      END
   END clk1
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER MET4 ;
         RECT  178.48 975.2 179.04 976.68 ;
      END
   END dout1[0]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER MET4 ;
         RECT  212.52 975.2 213.08 976.68 ;
      END
   END dout1[1]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER MET4 ;
         RECT  246.56 975.2 247.12 976.68 ;
      END
   END dout1[2]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER MET4 ;
         RECT  278.76 975.2 279.32 976.68 ;
      END
   END dout1[3]
   PIN dout1[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER MET4 ;
         RECT  312.8 975.2 313.36 976.68 ;
      END
   END dout1[4]
   PIN dout1[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER MET4 ;
         RECT  347.76 975.2 348.32 976.68 ;
      END
   END dout1[5]
   PIN dout1[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER MET4 ;
         RECT  381.8 975.2 382.36 976.68 ;
      END
   END dout1[6]
   PIN dout1[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER MET4 ;
         RECT  415.84 975.2 416.4 976.68 ;
      END
   END dout1[7]
   PIN dout1[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER MET4 ;
         RECT  448.04 975.2 448.6 976.68 ;
      END
   END dout1[8]
   PIN dout1[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER MET4 ;
         RECT  482.08 975.2 482.64 976.68 ;
      END
   END dout1[9]
   PIN dout1[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER MET4 ;
         RECT  517.04 975.2 517.6 976.68 ;
      END
   END dout1[10]
   PIN dout1[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER MET4 ;
         RECT  551.08 975.2 551.64 976.68 ;
      END
   END dout1[11]
   PIN dout1[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER MET4 ;
         RECT  585.12 975.2 585.68 976.68 ;
      END
   END dout1[12]
   PIN dout1[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER MET4 ;
         RECT  617.32 975.2 617.88 976.68 ;
      END
   END dout1[13]
   PIN dout1[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER MET4 ;
         RECT  651.36 975.2 651.92 976.68 ;
      END
   END dout1[14]
   PIN dout1[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER MET4 ;
         RECT  686.32 975.2 686.88 976.68 ;
      END
   END dout1[15]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER MET4 ;
         RECT  530.84 0.0 531.4 976.68 ;
         LAYER MET4 ;
         RECT  823.4 0.0 823.96 976.68 ;
         LAYER MET3 ;
         RECT  0.0 792.12 899.4 792.68 ;
         LAYER MET3 ;
         RECT  0.0 928.28 899.4 928.84 ;
         LAYER MET3 ;
         RECT  821.56 54.28 899.4 54.84 ;
         LAYER MET3 ;
         RECT  755.32 863.88 899.4 864.44 ;
         LAYER MET4 ;
         RECT  205.16 14.72 205.72 976.68 ;
         LAYER MET4 ;
         RECT  379.96 0.0 380.52 976.68 ;
         LAYER MET3 ;
         RECT  0.0 190.44 160.64 191.0 ;
         LAYER MET3 ;
         RECT  0.0 959.56 766.0 960.12 ;
         LAYER MET4 ;
         RECT  852.84 0.0 853.4 976.68 ;
         LAYER MET3 ;
         RECT  0.0 76.36 815.68 76.92 ;
         LAYER MET4 ;
         RECT  348.68 20.24 349.24 976.68 ;
         LAYER MET4 ;
         RECT  381.8 0.0 382.36 9.76 ;
         LAYER MET3 ;
         RECT  780.16 194.12 899.4 194.68 ;
         LAYER MET3 ;
         RECT  0.0 343.16 899.4 343.72 ;
         LAYER MET3 ;
         RECT  716.68 396.52 899.4 397.08 ;
         LAYER MET3 ;
         RECT  405.72 2.76 899.4 3.32 ;
         LAYER MET4 ;
         RECT  109.48 0.0 110.04 976.68 ;
         LAYER MET3 ;
         RECT  780.16 243.8 899.4 244.36 ;
         LAYER MET3 ;
         RECT  0.0 48.76 185.48 49.32 ;
         LAYER MET3 ;
         RECT  0.0 280.6 117.4 281.16 ;
         LAYER MET3 ;
         RECT  716.68 446.2 899.4 446.76 ;
         LAYER MET3 ;
         RECT  0.0 735.08 899.4 735.64 ;
         LAYER MET4 ;
         RECT  59.8 0.0 60.36 976.68 ;
         LAYER MET4 ;
         RECT  243.8 6.44 244.36 976.68 ;
         LAYER MET4 ;
         RECT  554.76 0.0 555.32 976.68 ;
         LAYER MET4 ;
         RECT  792.12 0.0 792.68 976.68 ;
         LAYER MET3 ;
         RECT  0.0 797.64 899.4 798.2 ;
         LAYER MET3 ;
         RECT  0.0 483.0 899.4 483.56 ;
         LAYER MET3 ;
         RECT  0.0 98.44 117.4 99.0 ;
         LAYER MET3 ;
         RECT  721.28 931.96 899.4 932.52 ;
         LAYER MET4 ;
         RECT  746.12 0.0 746.68 976.68 ;
         LAYER MET4 ;
         RECT  678.04 0.0 678.6 976.68 ;
         LAYER MET3 ;
         RECT  0.0 269.56 117.4 270.12 ;
         LAYER MET3 ;
         RECT  755.32 315.56 899.4 316.12 ;
         LAYER MET4 ;
         RECT  501.4 0.0 501.96 976.68 ;
         LAYER MET4 ;
         RECT  271.4 0.0 271.96 5.16 ;
         LAYER MET3 ;
         RECT  0.0 306.36 899.4 306.92 ;
         LAYER MET3 ;
         RECT  733.24 317.4 899.4 317.96 ;
         LAYER MET3 ;
         RECT  0.0 451.72 899.4 452.28 ;
         LAYER MET3 ;
         RECT  0.0 931.96 185.48 932.52 ;
         LAYER MET4 ;
         RECT  431.48 0.0 432.04 976.68 ;
         LAYER MET3 ;
         RECT  0.0 459.08 177.2 459.64 ;
         LAYER MET3 ;
         RECT  0.0 639.4 142.24 639.96 ;
         LAYER MET3 ;
         RECT  0.0 760.84 899.4 761.4 ;
         LAYER MET4 ;
         RECT  6.44 0.0 7.0 976.68 ;
         LAYER MET4 ;
         RECT  506.92 0.0 507.48 976.68 ;
         LAYER MET4 ;
         RECT  862.04 0.0 862.6 959.2 ;
         LAYER MET3 ;
         RECT  0.0 720.36 177.2 720.92 ;
         LAYER MET4 ;
         RECT  799.48 0.0 800.04 976.68 ;
         LAYER MET4 ;
         RECT  492.2 0.0 492.76 976.68 ;
         LAYER MET4 ;
         RECT  819.72 46.0 820.28 976.68 ;
         LAYER MET3 ;
         RECT  0.0 348.68 899.4 349.24 ;
         LAYER MET4 ;
         RECT  451.72 0.0 452.28 976.68 ;
         LAYER MET4 ;
         RECT  271.4 16.56 271.96 976.68 ;
         LAYER MET4 ;
         RECT  116.84 0.0 117.4 976.68 ;
         LAYER MET3 ;
         RECT  0.0 970.6 752.2 971.16 ;
         LAYER MET3 ;
         RECT  0.0 365.24 142.24 365.8 ;
         LAYER MET3 ;
         RECT  0.0 729.56 899.4 730.12 ;
         LAYER MET4 ;
         RECT  626.52 0.0 627.08 976.68 ;
         LAYER MET4 ;
         RECT  663.32 0.0 663.88 976.68 ;
         LAYER MET4 ;
         RECT  692.76 0.0 693.32 976.68 ;
         LAYER MET3 ;
         RECT  716.68 832.6 899.4 833.16 ;
         LAYER MET4 ;
         RECT  332.12 0.0 332.68 976.68 ;
         LAYER MET3 ;
         RECT  0.0 89.24 804.64 89.8 ;
         LAYER MET3 ;
         RECT  0.0 319.24 77.84 319.8 ;
         LAYER MET3 ;
         RECT  755.32 788.44 899.4 789.0 ;
         LAYER MET3 ;
         RECT  0.0 538.2 162.48 538.76 ;
         LAYER MET3 ;
         RECT  0.0 591.56 899.4 592.12 ;
         LAYER MET4 ;
         RECT  495.88 0.0 496.44 976.68 ;
         LAYER MET4 ;
         RECT  720.36 0.0 720.92 976.68 ;
         LAYER MET3 ;
         RECT  780.16 183.08 899.4 183.64 ;
         LAYER MET3 ;
         RECT  0.0 523.48 899.4 524.04 ;
         LAYER MET4 ;
         RECT  142.6 0.0 143.16 976.68 ;
         LAYER MET3 ;
         RECT  0.0 768.2 899.4 768.76 ;
         LAYER MET4 ;
         RECT  203.32 0.0 203.88 976.68 ;
         LAYER MET4 ;
         RECT  315.56 20.24 316.12 976.68 ;
         LAYER MET4 ;
         RECT  808.68 0.0 809.24 976.68 ;
         LAYER MET4 ;
         RECT  341.32 0.0 341.88 976.68 ;
         LAYER MET4 ;
         RECT  387.32 12.88 387.88 976.68 ;
         LAYER MET3 ;
         RECT  0.0 593.4 899.4 593.96 ;
         LAYER MET3 ;
         RECT  716.68 148.12 899.4 148.68 ;
         LAYER MET3 ;
         RECT  0.0 400.2 899.4 400.76 ;
         LAYER MET3 ;
         RECT  809.6 933.8 899.4 934.36 ;
         LAYER MET4 ;
         RECT  460.92 0.0 461.48 976.68 ;
         LAYER MET3 ;
         RECT  0.0 586.04 899.4 586.6 ;
         LAYER MET3 ;
         RECT  0.0 293.48 73.24 294.04 ;
         LAYER MET4 ;
         RECT  311.88 0.0 312.44 976.68 ;
         LAYER MET3 ;
         RECT  0.0 391.0 142.24 391.56 ;
         LAYER MET3 ;
         RECT  0.0 322.92 177.2 323.48 ;
         LAYER MET4 ;
         RECT  78.2 0.0 78.76 976.68 ;
         LAYER MET3 ;
         RECT  0.0 23.0 121.08 23.56 ;
         LAYER MET3 ;
         RECT  0.0 173.88 177.2 174.44 ;
         LAYER MET3 ;
         RECT  0.0 628.36 899.4 628.92 ;
         LAYER MET4 ;
         RECT  4.6 0.0 5.16 976.68 ;
         LAYER MET3 ;
         RECT  0.0 679.88 899.4 680.44 ;
         LAYER MET4 ;
         RECT  105.8 0.0 106.36 976.68 ;
         LAYER MET3 ;
         RECT  0.0 808.68 899.4 809.24 ;
         LAYER MET4 ;
         RECT  641.24 0.0 641.8 976.68 ;
         LAYER MET3 ;
         RECT  0.0 448.04 899.4 448.6 ;
         LAYER MET4 ;
         RECT  895.16 0.0 895.72 976.68 ;
         LAYER MET3 ;
         RECT  0.0 948.52 899.4 949.08 ;
         LAYER MET3 ;
         RECT  0.0 118.68 117.4 119.24 ;
         LAYER MET4 ;
         RECT  133.4 0.0 133.96 976.68 ;
         LAYER MET3 ;
         RECT  0.0 966.92 899.4 967.48 ;
         LAYER MET3 ;
         RECT  716.68 819.72 899.4 820.28 ;
         LAYER MET3 ;
         RECT  0.0 339.48 160.64 340.04 ;
         LAYER MET4 ;
         RECT  455.4 0.0 455.96 976.68 ;
         LAYER MET4 ;
         RECT  199.64 0.0 200.2 976.68 ;
         LAYER MET4 ;
         RECT  718.52 0.0 719.08 976.68 ;
         LAYER MET3 ;
         RECT  780.16 210.68 899.4 211.24 ;
         LAYER MET4 ;
         RECT  57.96 0.0 58.52 976.68 ;
         LAYER MET3 ;
         RECT  0.0 582.36 899.4 582.92 ;
         LAYER MET3 ;
         RECT  733.24 289.8 899.4 290.36 ;
         LAYER MET3 ;
         RECT  0.0 203.32 117.4 203.88 ;
         LAYER MET4 ;
         RECT  83.72 0.0 84.28 976.68 ;
         LAYER MET4 ;
         RECT  619.16 0.0 619.72 17.12 ;
         LAYER MET3 ;
         RECT  0.0 906.2 882.84 906.76 ;
         LAYER MET4 ;
         RECT  155.48 0.0 156.04 5.16 ;
         LAYER MET3 ;
         RECT  0.0 687.24 899.4 687.8 ;
         LAYER MET4 ;
         RECT  541.88 0.0 542.44 976.68 ;
         LAYER MET4 ;
         RECT  438.84 0.0 439.4 976.68 ;
         LAYER MET3 ;
         RECT  0.0 775.56 899.4 776.12 ;
         LAYER MET3 ;
         RECT  0.0 621.0 177.2 621.56 ;
         LAYER MET3 ;
         RECT  0.0 828.92 899.4 829.48 ;
         LAYER MET3 ;
         RECT  0.0 904.36 899.4 904.92 ;
         LAYER MET4 ;
         RECT  15.64 0.0 16.2 976.68 ;
         LAYER MET3 ;
         RECT  0.0 663.32 160.64 663.88 ;
         LAYER MET3 ;
         RECT  0.0 411.24 899.4 411.8 ;
         LAYER MET4 ;
         RECT  232.76 0.0 233.32 976.68 ;
         LAYER MET4 ;
         RECT  300.84 0.0 301.4 976.68 ;
         LAYER MET4 ;
         RECT  475.64 0.0 476.2 976.68 ;
         LAYER MET4 ;
         RECT  740.6 0.0 741.16 976.68 ;
         LAYER MET4 ;
         RECT  102.12 0.0 102.68 976.68 ;
         LAYER MET4 ;
         RECT  289.8 0.0 290.36 976.68 ;
         LAYER MET4 ;
         RECT  409.4 0.0 409.96 976.68 ;
         LAYER MET4 ;
         RECT  797.64 0.0 798.2 976.68 ;
         LAYER MET3 ;
         RECT  0.0 398.36 899.4 398.92 ;
         LAYER MET4 ;
         RECT  654.12 0.0 654.68 9.76 ;
         LAYER MET3 ;
         RECT  0.0 333.96 177.2 334.52 ;
         LAYER MET3 ;
         RECT  0.0 356.04 899.4 356.6 ;
         LAYER MET3 ;
         RECT  0.0 28.52 30.92 29.08 ;
         LAYER MET3 ;
         RECT  0.0 933.8 739.32 934.36 ;
         LAYER MET3 ;
         RECT  0.0 852.84 899.4 853.4 ;
         LAYER MET4 ;
         RECT  619.16 20.24 619.72 976.68 ;
         LAYER MET4 ;
         RECT  549.24 0.0 549.8 976.68 ;
         LAYER MET3 ;
         RECT  821.56 63.48 899.4 64.04 ;
         LAYER MET3 ;
         RECT  0.0 525.32 899.4 525.88 ;
         LAYER MET3 ;
         RECT  733.24 762.68 899.4 763.24 ;
         LAYER MET3 ;
         RECT  716.68 297.16 899.4 297.72 ;
         LAYER MET3 ;
         RECT  0.0 968.76 899.4 969.32 ;
         LAYER MET4 ;
         RECT  184.92 0.0 185.48 976.68 ;
         LAYER MET3 ;
         RECT  0.0 102.12 899.4 102.68 ;
         LAYER MET3 ;
         RECT  0.0 880.44 899.4 881.0 ;
         LAYER MET3 ;
         RECT  0.0 793.96 899.4 794.52 ;
         LAYER MET3 ;
         RECT  731.4 740.6 899.4 741.16 ;
         LAYER MET3 ;
         RECT  91.08 24.84 899.4 25.4 ;
         LAYER MET4 ;
         RECT  337.64 18.4 338.2 976.68 ;
         LAYER MET4 ;
         RECT  420.44 0.0 421.0 976.68 ;
         LAYER MET3 ;
         RECT  0.0 192.28 100.84 192.84 ;
         LAYER MET3 ;
         RECT  733.24 516.12 899.4 516.68 ;
         LAYER MET3 ;
         RECT  755.32 365.24 899.4 365.8 ;
         LAYER MET3 ;
         RECT  780.16 133.4 899.4 133.96 ;
         LAYER MET3 ;
         RECT  0.0 930.12 808.32 930.68 ;
         LAYER MET3 ;
         RECT  0.0 414.92 142.24 415.48 ;
         LAYER MET3 ;
         RECT  0.0 289.8 160.64 290.36 ;
         LAYER MET3 ;
         RECT  0.0 703.8 899.4 704.36 ;
         LAYER MET3 ;
         RECT  0.0 197.8 117.4 198.36 ;
         LAYER MET3 ;
         RECT  780.16 278.76 899.4 279.32 ;
         LAYER MET3 ;
         RECT  0.0 372.6 177.2 373.16 ;
         LAYER MET3 ;
         RECT  780.16 286.12 899.4 286.68 ;
         LAYER MET3 ;
         RECT  0.0 367.08 160.64 367.64 ;
         LAYER MET3 ;
         RECT  0.0 740.6 162.48 741.16 ;
         LAYER MET4 ;
         RECT  639.4 0.0 639.96 976.68 ;
         LAYER MET3 ;
         RECT  0.0 913.56 158.8 914.12 ;
         LAYER MET4 ;
         RECT  711.16 0.0 711.72 976.68 ;
         LAYER MET3 ;
         RECT  739.68 908.04 899.4 908.6 ;
         LAYER MET4 ;
         RECT  569.48 0.0 570.04 976.68 ;
         LAYER MET3 ;
         RECT  0.0 816.04 899.4 816.6 ;
         LAYER MET4 ;
         RECT  247.48 20.24 248.04 976.68 ;
         LAYER MET4 ;
         RECT  529.0 0.0 529.56 976.68 ;
         LAYER MET3 ;
         RECT  0.0 860.2 881.0 860.76 ;
         LAYER MET4 ;
         RECT  672.52 0.0 673.08 976.68 ;
         LAYER MET3 ;
         RECT  755.32 814.2 899.4 814.76 ;
         LAYER MET3 ;
         RECT  0.0 437.0 899.4 437.56 ;
         LAYER MET3 ;
         RECT  780.16 205.16 899.4 205.72 ;
         LAYER MET4 ;
         RECT  422.28 0.0 422.84 976.68 ;
         LAYER MET3 ;
         RECT  0.0 527.16 899.4 527.72 ;
         LAYER MET4 ;
         RECT  275.08 0.0 275.64 976.68 ;
         LAYER MET3 ;
         RECT  0.0 635.72 899.4 636.28 ;
         LAYER MET3 ;
         RECT  0.0 179.4 117.4 179.96 ;
         LAYER MET4 ;
         RECT  863.88 0.0 864.44 976.68 ;
         LAYER MET3 ;
         RECT  0.0 409.4 177.2 409.96 ;
         LAYER MET3 ;
         RECT  0.0 917.24 752.2 917.8 ;
         LAYER MET3 ;
         RECT  405.72 6.44 899.4 7.0 ;
         LAYER MET3 ;
         RECT  733.24 416.76 899.4 417.32 ;
         LAYER MET3 ;
         RECT  0.0 543.72 899.4 544.28 ;
         LAYER MET4 ;
         RECT  76.36 0.0 76.92 976.68 ;
         LAYER MET4 ;
         RECT  464.6 0.0 465.16 976.68 ;
         LAYER MET4 ;
         RECT  510.6 0.0 511.16 976.68 ;
         LAYER MET3 ;
         RECT  0.0 164.68 899.4 165.24 ;
         LAYER MET3 ;
         RECT  0.0 516.12 160.64 516.68 ;
         LAYER MET4 ;
         RECT  768.2 0.0 768.76 976.68 ;
         LAYER MET4 ;
         RECT  643.08 0.0 643.64 976.68 ;
         LAYER MET4 ;
         RECT  565.8 0.0 566.36 976.68 ;
         LAYER MET4 ;
         RECT  617.32 0.0 617.88 962.88 ;
         LAYER MET3 ;
         RECT  0.0 464.6 142.24 465.16 ;
         LAYER MET3 ;
         RECT  0.0 85.56 177.2 86.12 ;
         LAYER MET3 ;
         RECT  0.0 554.76 899.4 555.32 ;
         LAYER MET3 ;
         RECT  0.0 19.32 179.04 19.88 ;
         LAYER MET3 ;
         RECT  94.76 304.52 899.4 305.08 ;
         LAYER MET4 ;
         RECT  591.56 0.0 592.12 976.68 ;
         LAYER MET3 ;
         RECT  0.0 832.6 177.2 833.16 ;
         LAYER MET4 ;
         RECT  151.8 0.0 152.36 976.68 ;
         LAYER MET3 ;
         RECT  797.64 192.28 899.4 192.84 ;
         LAYER MET3 ;
         RECT  780.16 170.2 899.4 170.76 ;
         LAYER MET3 ;
         RECT  0.0 685.4 899.4 685.96 ;
         LAYER MET3 ;
         RECT  0.0 661.48 899.4 662.04 ;
         LAYER MET3 ;
         RECT  0.0 2.76 89.8 3.32 ;
         LAYER MET3 ;
         RECT  716.68 621.0 899.4 621.56 ;
         LAYER MET3 ;
         RECT  0.0 839.96 160.64 840.52 ;
         LAYER MET3 ;
         RECT  0.0 444.36 899.4 444.92 ;
         LAYER MET3 ;
         RECT  0.0 950.36 856.16 950.92 ;
         LAYER MET4 ;
         RECT  413.08 0.0 413.64 976.68 ;
         LAYER MET3 ;
         RECT  0.0 838.12 142.24 838.68 ;
         LAYER MET3 ;
         RECT  0.0 61.64 89.8 62.2 ;
         LAYER MET3 ;
         RECT  0.0 547.4 899.4 547.96 ;
         LAYER MET4 ;
         RECT  536.36 0.0 536.92 976.68 ;
         LAYER MET4 ;
         RECT  356.04 0.0 356.6 976.68 ;
         LAYER MET4 ;
         RECT  604.44 0.0 605.0 976.68 ;
         LAYER MET3 ;
         RECT  0.0 499.56 899.4 500.12 ;
         LAYER MET3 ;
         RECT  0.0 619.16 899.4 619.72 ;
         LAYER MET4 ;
         RECT  650.44 0.0 651.0 962.88 ;
         LAYER MET4 ;
         RECT  374.44 0.0 375.0 976.68 ;
         LAYER MET3 ;
         RECT  797.64 291.64 899.4 292.2 ;
         LAYER MET3 ;
         RECT  0.0 142.6 100.84 143.16 ;
         LAYER MET3 ;
         RECT  0.0 416.76 160.64 417.32 ;
         LAYER MET3 ;
         RECT  733.24 69.0 899.4 69.56 ;
         LAYER MET3 ;
         RECT  0.0 131.56 117.4 132.12 ;
         LAYER MET3 ;
         RECT  0.0 291.64 80.6 292.2 ;
         LAYER MET3 ;
         RECT  733.24 839.96 899.4 840.52 ;
         LAYER MET3 ;
         RECT  780.16 94.76 899.4 95.32 ;
         LAYER MET3 ;
         RECT  755.32 838.12 899.4 838.68 ;
         LAYER MET4 ;
         RECT  287.96 14.72 288.52 976.68 ;
         LAYER MET4 ;
         RECT  731.4 0.0 731.96 976.68 ;
         LAYER MET3 ;
         RECT  780.16 184.92 899.4 185.48 ;
         LAYER MET3 ;
         RECT  0.0 935.64 899.4 936.2 ;
         LAYER MET4 ;
         RECT  394.68 0.0 395.24 976.68 ;
         LAYER MET3 ;
         RECT  0.0 59.8 899.4 60.36 ;
         LAYER MET4 ;
         RECT  777.4 0.0 777.96 976.68 ;
         LAYER MET3 ;
         RECT  0.0 510.6 899.4 511.16 ;
         LAYER MET3 ;
         RECT  0.0 654.12 899.4 654.68 ;
         LAYER MET3 ;
         RECT  780.16 247.48 899.4 248.04 ;
         LAYER MET3 ;
         RECT  0.0 560.28 899.4 560.84 ;
         LAYER MET4 ;
         RECT  251.16 0.0 251.72 976.68 ;
         LAYER MET3 ;
         RECT  0.0 275.08 899.4 275.64 ;
         LAYER MET3 ;
         RECT  0.0 389.16 160.64 389.72 ;
         LAYER MET3 ;
         RECT  0.0 556.6 899.4 557.16 ;
         LAYER MET3 ;
         RECT  892.4 854.68 899.4 855.24 ;
         LAYER MET4 ;
         RECT  35.88 0.0 36.44 976.68 ;
         LAYER MET3 ;
         RECT  0.0 718.52 899.4 719.08 ;
         LAYER MET3 ;
         RECT  0.0 891.48 899.4 892.04 ;
         LAYER MET3 ;
         RECT  0.0 937.48 899.4 938.04 ;
         LAYER MET4 ;
         RECT  725.88 0.0 726.44 976.68 ;
         LAYER MET3 ;
         RECT  0.0 181.24 117.4 181.8 ;
         LAYER MET3 ;
         RECT  0.0 10.12 5.16 10.68 ;
         LAYER MET4 ;
         RECT  221.72 0.0 222.28 5.16 ;
         LAYER MET3 ;
         RECT  0.0 519.8 899.4 520.36 ;
         LAYER MET3 ;
         RECT  0.0 194.12 117.4 194.68 ;
         LAYER MET3 ;
         RECT  0.0 713.0 160.64 713.56 ;
         LAYER MET3 ;
         RECT  0.0 188.6 899.4 189.16 ;
         LAYER MET3 ;
         RECT  716.68 310.04 899.4 310.6 ;
         LAYER MET3 ;
         RECT  0.0 271.4 117.4 271.96 ;
         LAYER MET4 ;
         RECT  615.48 0.0 616.04 976.68 ;
         LAYER MET4 ;
         RECT  435.16 0.0 435.72 976.68 ;
         LAYER MET3 ;
         RECT  0.0 952.2 899.4 952.76 ;
         LAYER MET3 ;
         RECT  780.16 120.52 899.4 121.08 ;
         LAYER MET3 ;
         RECT  0.0 57.96 87.96 58.52 ;
         LAYER MET3 ;
         RECT  0.0 630.2 899.4 630.76 ;
         LAYER MET3 ;
         RECT  780.16 168.36 899.4 168.92 ;
         LAYER MET3 ;
         RECT  0.0 843.64 899.4 844.2 ;
         LAYER MET3 ;
         RECT  0.0 911.72 160.64 912.28 ;
         LAYER MET4 ;
         RECT  519.8 0.0 520.36 976.68 ;
         LAYER MET4 ;
         RECT  416.76 0.0 417.32 13.44 ;
         LAYER MET4 ;
         RECT  278.76 0.0 279.32 962.88 ;
         LAYER MET4 ;
         RECT  575.0 0.0 575.56 976.68 ;
         LAYER MET3 ;
         RECT  0.0 394.68 899.4 395.24 ;
         LAYER MET3 ;
         RECT  771.88 970.6 899.4 971.16 ;
         LAYER MET4 ;
         RECT  144.44 6.44 145.0 976.68 ;
         LAYER MET3 ;
         RECT  0.0 954.04 849.72 954.6 ;
         LAYER MET4 ;
         RECT  28.52 0.0 29.08 976.68 ;
         LAYER MET4 ;
         RECT  229.08 0.0 229.64 976.68 ;
         LAYER MET4 ;
         RECT  234.6 0.0 235.16 976.68 ;
         LAYER MET3 ;
         RECT  0.0 541.88 899.4 542.44 ;
         LAYER MET4 ;
         RECT  701.96 0.0 702.52 976.68 ;
         LAYER MET4 ;
         RECT  195.96 0.0 196.52 976.68 ;
         LAYER MET3 ;
         RECT  83.72 308.2 899.4 308.76 ;
         LAYER MET3 ;
         RECT  716.68 608.12 899.4 608.68 ;
         LAYER MET3 ;
         RECT  0.0 595.24 177.2 595.8 ;
         LAYER MET4 ;
         RECT  256.68 0.0 257.24 976.68 ;
         LAYER MET3 ;
         RECT  0.0 939.32 899.4 939.88 ;
         LAYER MET3 ;
         RECT  0.0 909.88 881.0 910.44 ;
         LAYER MET4 ;
         RECT  749.8 0.0 750.36 976.68 ;
         LAYER MET4 ;
         RECT  449.88 20.24 450.44 976.68 ;
         LAYER MET3 ;
         RECT  0.0 381.8 899.4 382.36 ;
         LAYER MET3 ;
         RECT  0.0 457.24 899.4 457.8 ;
         LAYER MET3 ;
         RECT  97.52 328.44 899.4 329.0 ;
         LAYER MET3 ;
         RECT  0.0 563.96 142.24 564.52 ;
         LAYER MET3 ;
         RECT  733.24 663.32 899.4 663.88 ;
         LAYER MET3 ;
         RECT  755.32 738.76 899.4 739.32 ;
         LAYER MET4 ;
         RECT  264.04 0.0 264.6 976.68 ;
         LAYER MET4 ;
         RECT  497.72 0.0 498.28 976.68 ;
         LAYER MET3 ;
         RECT  0.0 177.56 899.4 178.12 ;
         LAYER MET3 ;
         RECT  0.0 694.6 899.4 695.16 ;
         LAYER MET3 ;
         RECT  0.0 420.44 899.4 421.0 ;
         LAYER MET3 ;
         RECT  0.0 427.8 899.4 428.36 ;
         LAYER MET3 ;
         RECT  0.0 225.4 899.4 225.96 ;
         LAYER MET3 ;
         RECT  0.0 757.16 177.2 757.72 ;
         LAYER MET4 ;
         RECT  700.12 0.0 700.68 976.68 ;
         LAYER MET4 ;
         RECT  865.72 0.0 866.28 976.68 ;
         LAYER MET3 ;
         RECT  0.0 341.32 80.6 341.88 ;
         LAYER MET3 ;
         RECT  0.0 862.04 160.64 862.6 ;
         LAYER MET3 ;
         RECT  0.0 957.72 864.44 958.28 ;
         LAYER MET3 ;
         RECT  0.0 644.92 899.4 645.48 ;
         LAYER MET4 ;
         RECT  267.72 0.0 268.28 976.68 ;
         LAYER MET3 ;
         RECT  733.24 911.72 899.4 912.28 ;
         LAYER MET4 ;
         RECT  280.6 0.0 281.16 11.6 ;
         LAYER MET4 ;
         RECT  571.32 0.0 571.88 976.68 ;
         LAYER MET4 ;
         RECT  560.28 0.0 560.84 976.68 ;
         LAYER MET3 ;
         RECT  0.0 781.08 899.4 781.64 ;
         LAYER MET3 ;
         RECT  797.64 216.2 899.4 216.76 ;
         LAYER MET3 ;
         RECT  0.0 148.12 177.2 148.68 ;
         LAYER MET3 ;
         RECT  0.0 247.48 117.4 248.04 ;
         LAYER MET4 ;
         RECT  37.72 0.0 38.28 976.68 ;
         LAYER MET3 ;
         RECT  821.56 61.64 899.4 62.2 ;
         LAYER MET4 ;
         RECT  378.12 0.0 378.68 976.68 ;
         LAYER MET3 ;
         RECT  0.0 265.88 100.84 266.44 ;
         LAYER MET4 ;
         RECT  91.08 0.0 91.64 976.68 ;
         LAYER MET3 ;
         RECT  0.0 267.72 117.4 268.28 ;
         LAYER MET3 ;
         RECT  0.0 744.28 899.4 744.84 ;
         LAYER MET4 ;
         RECT  538.2 0.0 538.76 976.68 ;
         LAYER MET4 ;
         RECT  795.8 0.0 796.36 976.68 ;
         LAYER MET4 ;
         RECT  816.04 0.0 816.6 976.68 ;
         LAYER MET4 ;
         RECT  606.28 0.0 606.84 976.68 ;
         LAYER MET4 ;
         RECT  885.96 0.0 886.52 976.68 ;
         LAYER MET3 ;
         RECT  755.32 887.8 899.4 888.36 ;
         LAYER MET3 ;
         RECT  0.0 849.16 899.4 849.72 ;
         LAYER MET3 ;
         RECT  0.0 606.28 899.4 606.84 ;
         LAYER MET4 ;
         RECT  21.16 0.0 21.72 976.68 ;
         LAYER MET4 ;
         RECT  39.56 0.0 40.12 976.68 ;
         LAYER MET4 ;
         RECT  291.64 0.0 292.2 976.68 ;
         LAYER MET4 ;
         RECT  403.88 0.0 404.44 5.16 ;
         LAYER MET4 ;
         RECT  512.44 0.0 513.0 976.68 ;
         LAYER MET3 ;
         RECT  755.32 540.04 899.4 540.6 ;
         LAYER MET3 ;
         RECT  0.0 100.28 7.0 100.84 ;
         LAYER MET3 ;
         RECT  0.0 900.68 899.4 901.24 ;
         LAYER MET3 ;
         RECT  83.72 324.76 899.4 325.32 ;
         LAYER MET3 ;
         RECT  0.0 144.44 899.4 145.0 ;
         LAYER MET3 ;
         RECT  755.32 464.6 899.4 465.16 ;
         LAYER MET3 ;
         RECT  0.0 648.6 899.4 649.16 ;
         LAYER MET3 ;
         RECT  0.0 497.72 899.4 498.28 ;
         LAYER MET3 ;
         RECT  716.68 173.88 899.4 174.44 ;
         LAYER MET4 ;
         RECT  521.64 0.0 522.2 976.68 ;
         LAYER MET4 ;
         RECT  757.16 0.0 757.72 976.68 ;
         LAYER MET3 ;
         RECT  0.0 696.44 899.4 697.0 ;
         LAYER MET3 ;
         RECT  0.0 874.92 899.4 875.48 ;
         LAYER MET4 ;
         RECT  339.48 0.0 340.04 976.68 ;
         LAYER MET4 ;
         RECT  611.8 0.0 612.36 976.68 ;
         LAYER MET3 ;
         RECT  0.0 766.36 899.4 766.92 ;
         LAYER MET4 ;
         RECT  418.6 0.0 419.16 976.68 ;
         LAYER MET3 ;
         RECT  0.0 786.6 899.4 787.16 ;
         LAYER MET3 ;
         RECT  780.16 172.04 899.4 172.6 ;
         LAYER MET3 ;
         RECT  0.0 512.44 899.4 513.0 ;
         LAYER MET3 ;
         RECT  0.0 284.28 117.4 284.84 ;
         LAYER MET4 ;
         RECT  810.52 0.0 811.08 976.68 ;
         LAYER MET4 ;
         RECT  241.96 0.0 242.52 976.68 ;
         LAYER MET4 ;
         RECT  889.64 0.0 890.2 976.68 ;
         LAYER MET3 ;
         RECT  780.16 273.24 899.4 273.8 ;
         LAYER MET4 ;
         RECT  162.84 0.0 163.4 976.68 ;
         LAYER MET3 ;
         RECT  0.0 376.28 899.4 376.84 ;
         LAYER MET3 ;
         RECT  0.0 747.96 899.4 748.52 ;
         LAYER MET3 ;
         RECT  0.0 963.24 176.28 963.8 ;
         LAYER MET4 ;
         RECT  302.68 0.0 303.24 976.68 ;
         LAYER MET4 ;
         RECT  219.88 0.0 220.44 976.68 ;
         LAYER MET4 ;
         RECT  867.56 0.0 868.12 976.68 ;
         LAYER MET4 ;
         RECT  753.48 0.0 754.04 976.68 ;
         LAYER MET3 ;
         RECT  0.0 819.72 177.2 820.28 ;
         LAYER MET4 ;
         RECT  667.0 0.0 667.56 976.68 ;
         LAYER MET3 ;
         RECT  0.0 429.64 899.4 430.2 ;
         LAYER MET3 ;
         RECT  0.0 821.56 899.4 822.12 ;
         LAYER MET4 ;
         RECT  411.24 0.0 411.8 976.68 ;
         LAYER MET4 ;
         RECT  46.92 0.0 47.48 976.68 ;
         LAYER MET3 ;
         RECT  0.0 166.52 100.84 167.08 ;
         LAYER MET3 ;
         RECT  733.24 190.44 899.4 191.0 ;
         LAYER MET3 ;
         RECT  716.68 707.48 899.4 708.04 ;
         LAYER MET3 ;
         RECT  0.0 851.0 899.4 851.56 ;
         LAYER MET3 ;
         RECT  0.0 221.72 899.4 222.28 ;
         LAYER MET4 ;
         RECT  107.64 0.0 108.2 976.68 ;
         LAYER MET3 ;
         RECT  0.0 230.92 899.4 231.48 ;
         LAYER MET4 ;
         RECT  587.88 0.0 588.44 976.68 ;
         LAYER MET3 ;
         RECT  0.0 313.72 899.4 314.28 ;
         LAYER MET3 ;
         RECT  733.24 240.12 899.4 240.68 ;
         LAYER MET3 ;
         RECT  0.0 668.84 899.4 669.4 ;
         LAYER MET4 ;
         RECT  437.0 0.0 437.56 976.68 ;
         LAYER MET3 ;
         RECT  716.68 359.72 899.4 360.28 ;
         LAYER MET4 ;
         RECT  659.64 0.0 660.2 976.68 ;
         LAYER MET4 ;
         RECT  893.32 0.0 893.88 976.68 ;
         LAYER MET3 ;
         RECT  17.48 83.72 899.4 84.28 ;
         LAYER MET4 ;
         RECT  225.4 0.0 225.96 976.68 ;
         LAYER MET3 ;
         RECT  0.0 689.08 142.24 689.64 ;
         LAYER MET3 ;
         RECT  0.0 598.92 899.4 599.48 ;
         LAYER MET3 ;
         RECT  0.0 208.84 117.4 209.4 ;
         LAYER MET3 ;
         RECT  733.24 389.16 899.4 389.72 ;
         LAYER MET3 ;
         RECT  0.0 674.36 899.4 674.92 ;
         LAYER MET3 ;
         RECT  0.0 690.92 162.48 691.48 ;
         LAYER MET3 ;
         RECT  0.0 955.88 899.4 956.44 ;
         LAYER MET3 ;
         RECT  780.16 105.8 899.4 106.36 ;
         LAYER MET3 ;
         RECT  0.0 138.92 899.4 139.48 ;
         LAYER MET4 ;
         RECT  98.44 0.0 99.0 976.68 ;
         LAYER MET4 ;
         RECT  168.36 0.0 168.92 976.68 ;
         LAYER MET4 ;
         RECT  735.08 0.0 735.64 976.68 ;
         LAYER MET3 ;
         RECT  0.0 575.0 899.4 575.56 ;
         LAYER MET3 ;
         RECT  0.0 924.6 720.0 925.16 ;
         LAYER MET4 ;
         RECT  126.04 0.0 126.6 976.68 ;
         LAYER MET3 ;
         RECT  0.0 107.64 117.4 108.2 ;
         LAYER MET3 ;
         RECT  0.0 219.88 899.4 220.44 ;
         LAYER MET4 ;
         RECT  313.72 0.0 314.28 976.68 ;
         LAYER MET4 ;
         RECT  707.48 0.0 708.04 976.68 ;
         LAYER MET3 ;
         RECT  755.32 615.48 899.4 616.04 ;
         LAYER MET3 ;
         RECT  0.0 532.68 899.4 533.24 ;
         LAYER MET3 ;
         RECT  0.0 919.08 881.0 919.64 ;
         LAYER MET4 ;
         RECT  784.76 0.0 785.32 976.68 ;
         LAYER MET3 ;
         RECT  0.0 403.88 899.4 404.44 ;
         LAYER MET3 ;
         RECT  0.0 17.48 30.0 18.04 ;
         LAYER MET4 ;
         RECT  284.28 0.0 284.84 976.68 ;
         LAYER MET3 ;
         RECT  822.48 70.84 899.4 71.4 ;
         LAYER MET4 ;
         RECT  161.0 6.44 161.56 976.68 ;
         LAYER MET4 ;
         RECT  315.56 0.0 316.12 11.6 ;
         LAYER MET4 ;
         RECT  72.68 0.0 73.24 976.68 ;
         LAYER MET3 ;
         RECT  780.16 254.84 899.4 255.4 ;
         LAYER MET4 ;
         RECT  517.96 0.0 518.52 11.6 ;
         LAYER MET4 ;
         RECT  146.28 0.0 146.84 976.68 ;
         LAYER MET3 ;
         RECT  892.4 922.76 899.4 923.32 ;
         LAYER MET3 ;
         RECT  0.0 435.16 899.4 435.72 ;
         LAYER MET4 ;
         RECT  573.16 0.0 573.72 976.68 ;
         LAYER MET3 ;
         RECT  755.32 391.0 899.4 391.56 ;
         LAYER MET4 ;
         RECT  499.56 0.0 500.12 976.68 ;
         LAYER MET4 ;
         RECT  766.36 0.0 766.92 976.68 ;
         LAYER MET3 ;
         RECT  0.0 633.88 177.2 634.44 ;
         LAYER MET3 ;
         RECT  0.0 122.36 117.4 122.92 ;
         LAYER MET3 ;
         RECT  0.0 867.56 881.0 868.12 ;
         LAYER MET4 ;
         RECT  17.48 0.0 18.04 976.68 ;
         LAYER MET3 ;
         RECT  0.0 825.24 899.4 825.8 ;
         LAYER MET4 ;
         RECT  514.28 0.0 514.84 976.68 ;
         LAYER MET4 ;
         RECT  227.24 6.44 227.8 976.68 ;
         LAYER MET4 ;
         RECT  646.76 0.0 647.32 976.68 ;
         LAYER MET4 ;
         RECT  657.8 0.0 658.36 976.68 ;
         LAYER MET3 ;
         RECT  0.0 492.2 899.4 492.76 ;
         LAYER MET3 ;
         RECT  0.0 672.52 899.4 673.08 ;
         LAYER MET4 ;
         RECT  276.92 6.44 277.48 976.68 ;
         LAYER MET3 ;
         RECT  755.32 714.84 899.4 715.4 ;
         LAYER MET3 ;
         RECT  780.16 107.64 899.4 108.2 ;
         LAYER MET3 ;
         RECT  0.0 440.68 142.24 441.24 ;
         LAYER MET3 ;
         RECT  0.0 759.0 899.4 759.56 ;
         LAYER MET3 ;
         RECT  0.0 810.52 899.4 811.08 ;
         LAYER MET3 ;
         RECT  0.0 501.4 899.4 501.96 ;
         LAYER MET3 ;
         RECT  0.0 345.0 899.4 345.56 ;
         LAYER MET3 ;
         RECT  0.0 670.68 177.2 671.24 ;
         LAYER MET3 ;
         RECT  817.88 92.92 899.4 93.48 ;
         LAYER MET4 ;
         RECT  652.28 0.0 652.84 976.68 ;
         LAYER MET4 ;
         RECT  466.44 0.0 467.0 976.68 ;
         LAYER MET4 ;
         RECT  210.68 6.44 211.24 976.68 ;
         LAYER MET4 ;
         RECT  479.32 0.0 479.88 976.68 ;
         LAYER MET3 ;
         RECT  0.0 770.04 177.2 770.6 ;
         LAYER MET3 ;
         RECT  0.0 777.4 899.4 777.96 ;
         LAYER MET4 ;
         RECT  805.0 0.0 805.56 976.68 ;
         LAYER MET3 ;
         RECT  158.24 37.72 899.4 38.28 ;
         LAYER MET3 ;
         RECT  0.0 830.76 899.4 831.32 ;
         LAYER MET4 ;
         RECT  214.36 0.0 214.92 976.68 ;
         LAYER MET3 ;
         RECT  0.0 78.2 818.44 78.76 ;
         LAYER MET3 ;
         RECT  0.0 135.24 117.4 135.8 ;
         LAYER MET4 ;
         RECT  683.56 0.0 684.12 976.68 ;
         LAYER MET3 ;
         RECT  0.0 716.68 899.4 717.24 ;
         LAYER MET4 ;
         RECT  179.4 20.24 179.96 976.68 ;
         LAYER MET4 ;
         RECT  722.2 0.0 722.76 976.68 ;
         LAYER MET4 ;
         RECT  771.88 0.0 772.44 976.68 ;
         LAYER MET3 ;
         RECT  0.0 517.96 899.4 518.52 ;
         LAYER MET3 ;
         RECT  716.68 895.16 899.4 895.72 ;
         LAYER MET4 ;
         RECT  396.52 0.0 397.08 976.68 ;
         LAYER MET3 ;
         RECT  0.0 116.84 7.0 117.4 ;
         LAYER MET4 ;
         RECT  759.0 0.0 759.56 976.68 ;
         LAYER MET3 ;
         RECT  0.0 617.32 899.4 617.88 ;
         LAYER MET4 ;
         RECT  716.68 0.0 717.24 976.68 ;
         LAYER MET3 ;
         RECT  80.04 335.8 899.4 336.36 ;
         LAYER MET3 ;
         RECT  716.68 346.84 899.4 347.4 ;
         LAYER MET3 ;
         RECT  0.0 736.92 899.4 737.48 ;
         LAYER MET4 ;
         RECT  41.4 0.0 41.96 976.68 ;
         LAYER MET3 ;
         RECT  0.0 733.24 177.2 733.8 ;
         LAYER MET3 ;
         RECT  0.0 438.84 162.48 439.4 ;
         LAYER MET3 ;
         RECT  810.52 913.56 899.4 914.12 ;
         LAYER MET3 ;
         RECT  780.16 118.68 899.4 119.24 ;
         LAYER MET3 ;
         RECT  0.0 91.08 160.64 91.64 ;
         LAYER MET3 ;
         RECT  716.68 372.6 899.4 373.16 ;
         LAYER MET3 ;
         RECT  0.0 897.0 899.4 897.56 ;
         LAYER MET3 ;
         RECT  0.0 920.92 899.4 921.48 ;
         LAYER MET3 ;
         RECT  0.0 35.88 899.4 36.44 ;
         LAYER MET4 ;
         RECT  348.68 0.0 349.24 13.44 ;
         LAYER MET4 ;
         RECT  166.52 0.0 167.08 976.68 ;
         LAYER MET3 ;
         RECT  0.0 127.88 899.4 128.44 ;
         LAYER MET3 ;
         RECT  0.0 249.32 899.4 249.88 ;
         LAYER MET3 ;
         RECT  0.0 946.68 180.88 947.24 ;
         LAYER MET4 ;
         RECT  527.16 0.0 527.72 976.68 ;
         LAYER MET3 ;
         RECT  716.68 770.04 899.4 770.6 ;
         LAYER MET3 ;
         RECT  0.0 521.64 177.2 522.2 ;
         LAYER MET4 ;
         RECT  448.04 0.0 448.6 962.88 ;
         LAYER MET4 ;
         RECT  534.52 0.0 535.08 976.68 ;
         LAYER MET4 ;
         RECT  543.72 0.0 544.28 976.68 ;
         LAYER MET4 ;
         RECT  304.52 0.0 305.08 5.16 ;
         LAYER MET4 ;
         RECT  633.88 0.0 634.44 976.68 ;
         LAYER MET4 ;
         RECT  247.48 0.0 248.04 9.76 ;
         LAYER MET3 ;
         RECT  0.0 481.16 899.4 481.72 ;
         LAYER MET4 ;
         RECT  54.28 0.0 54.84 976.68 ;
         LAYER MET3 ;
         RECT  0.0 624.68 899.4 625.24 ;
         LAYER MET3 ;
         RECT  0.0 418.6 899.4 419.16 ;
         LAYER MET4 ;
         RECT  602.6 0.0 603.16 976.68 ;
         LAYER MET4 ;
         RECT  517.96 20.24 518.52 976.68 ;
         LAYER MET4 ;
         RECT  689.08 0.0 689.64 976.68 ;
         LAYER MET3 ;
         RECT  755.32 665.16 899.4 665.72 ;
         LAYER MET3 ;
         RECT  0.0 667.0 899.4 667.56 ;
         LAYER MET3 ;
         RECT  821.56 78.2 899.4 78.76 ;
         LAYER MET4 ;
         RECT  782.92 0.0 783.48 976.68 ;
         LAYER MET3 ;
         RECT  0.0 751.64 899.4 752.2 ;
         LAYER MET4 ;
         RECT  61.64 0.0 62.2 976.68 ;
         LAYER MET3 ;
         RECT  0.0 260.36 117.4 260.92 ;
         LAYER MET4 ;
         RECT  159.16 0.0 159.72 976.68 ;
         LAYER MET3 ;
         RECT  731.4 488.52 899.4 489.08 ;
         LAYER MET3 ;
         RECT  716.68 757.16 899.4 757.72 ;
         LAYER MET4 ;
         RECT  357.88 0.0 358.44 976.68 ;
         LAYER MET3 ;
         RECT  0.0 449.88 899.4 450.44 ;
         LAYER MET3 ;
         RECT  43.24 21.16 899.4 21.72 ;
         LAYER MET3 ;
         RECT  780.16 109.48 899.4 110.04 ;
         LAYER MET3 ;
         RECT  0.0 67.16 7.0 67.72 ;
         LAYER MET3 ;
         RECT  0.0 655.96 899.4 656.52 ;
         LAYER MET4 ;
         RECT  608.12 0.0 608.68 976.68 ;
         LAYER MET4 ;
         RECT  694.6 0.0 695.16 976.68 ;
         LAYER MET3 ;
         RECT  0.0 580.52 899.4 581.08 ;
         LAYER MET3 ;
         RECT  0.0 212.52 899.4 213.08 ;
         LAYER MET3 ;
         RECT  0.0 854.68 882.84 855.24 ;
         LAYER MET4 ;
         RECT  238.28 0.0 238.84 5.16 ;
         LAYER MET3 ;
         RECT  716.68 85.56 899.4 86.12 ;
         LAYER MET3 ;
         RECT  0.0 392.84 899.4 393.4 ;
         LAYER MET3 ;
         RECT  716.68 571.32 899.4 571.88 ;
         LAYER MET4 ;
         RECT  834.44 0.0 835.0 976.68 ;
         LAYER MET3 ;
         RECT  0.0 297.16 177.2 297.72 ;
         LAYER MET3 ;
         RECT  0.0 223.56 177.2 224.12 ;
         LAYER MET3 ;
         RECT  0.0 352.36 899.4 352.92 ;
         LAYER MET3 ;
         RECT  0.0 711.16 899.4 711.72 ;
         LAYER MET3 ;
         RECT  716.68 806.84 899.4 807.4 ;
         LAYER MET4 ;
         RECT  838.12 0.0 838.68 976.68 ;
         LAYER MET4 ;
         RECT  69.0 0.0 69.56 976.68 ;
         LAYER MET4 ;
         RECT  398.36 0.0 398.92 976.68 ;
         LAYER MET4 ;
         RECT  847.32 0.0 847.88 976.68 ;
         LAYER MET4 ;
         RECT  897.0 0.0 897.56 976.68 ;
         LAYER MET4 ;
         RECT  368.92 0.0 369.48 976.68 ;
         LAYER MET3 ;
         RECT  0.0 597.08 899.4 597.64 ;
         LAYER MET3 ;
         RECT  716.68 508.76 899.4 509.32 ;
         LAYER MET4 ;
         RECT  100.28 0.0 100.84 976.68 ;
         LAYER MET3 ;
         RECT  0.0 637.56 899.4 638.12 ;
         LAYER MET4 ;
         RECT  212.52 0.0 213.08 11.6 ;
         LAYER MET4 ;
         RECT  462.76 0.0 463.32 976.68 ;
         LAYER MET4 ;
         RECT  306.36 0.0 306.92 976.68 ;
         LAYER MET4 ;
         RECT  505.08 0.0 505.64 976.68 ;
         LAYER MET4 ;
         RECT  94.76 0.0 95.32 976.68 ;
         LAYER MET3 ;
         RECT  0.0 530.84 899.4 531.4 ;
         LAYER MET3 ;
         RECT  821.56 56.12 899.4 56.68 ;
         LAYER MET4 ;
         RECT  19.32 0.0 19.88 976.68 ;
         LAYER MET3 ;
         RECT  98.44 337.64 899.4 338.2 ;
         LAYER MET3 ;
         RECT  0.0 350.52 899.4 351.08 ;
         LAYER MET3 ;
         RECT  0.0 488.52 162.48 489.08 ;
         LAYER MET3 ;
         RECT  0.0 908.04 158.8 908.6 ;
         LAYER MET3 ;
         RECT  0.0 227.24 899.4 227.8 ;
         LAYER MET4 ;
         RECT  516.12 0.0 516.68 962.88 ;
         LAYER MET3 ;
         RECT  0.0 129.72 117.4 130.28 ;
         LAYER MET3 ;
         RECT  0.0 258.52 117.4 259.08 ;
         LAYER MET3 ;
         RECT  0.0 363.4 899.4 363.96 ;
         LAYER MET4 ;
         RECT  887.8 0.0 888.36 976.68 ;
         LAYER MET3 ;
         RECT  0.0 34.04 899.4 34.6 ;
         LAYER MET4 ;
         RECT  593.4 0.0 593.96 976.68 ;
         LAYER MET3 ;
         RECT  0.0 186.76 899.4 187.32 ;
         LAYER MET3 ;
         RECT  0.0 4.6 110.04 5.16 ;
         LAYER MET3 ;
         RECT  0.0 81.88 899.4 82.44 ;
         LAYER MET3 ;
         RECT  0.0 278.76 117.4 279.32 ;
         LAYER MET4 ;
         RECT  552.92 0.0 553.48 976.68 ;
         LAYER MET3 ;
         RECT  0.0 771.88 899.4 772.44 ;
         LAYER MET3 ;
         RECT  0.0 468.28 899.4 468.84 ;
         LAYER MET3 ;
         RECT  780.16 284.28 899.4 284.84 ;
         LAYER MET3 ;
         RECT  0.0 587.88 899.4 588.44 ;
         LAYER MET3 ;
         RECT  0.0 611.8 899.4 612.36 ;
         LAYER MET4 ;
         RECT  122.36 0.0 122.92 976.68 ;
         LAYER MET3 ;
         RECT  0.0 359.72 177.2 360.28 ;
         LAYER MET4 ;
         RECT  183.08 0.0 183.64 976.68 ;
         LAYER MET3 ;
         RECT  0.0 253.0 899.4 253.56 ;
         LAYER MET3 ;
         RECT  0.0 885.96 899.4 886.52 ;
         LAYER MET4 ;
         RECT  668.84 0.0 669.4 976.68 ;
         LAYER MET3 ;
         RECT  731.4 538.2 899.4 538.76 ;
         LAYER MET3 ;
         RECT  780.16 271.4 899.4 271.96 ;
         LAYER MET4 ;
         RECT  449.88 0.0 450.44 11.6 ;
         LAYER MET3 ;
         RECT  17.48 100.28 899.4 100.84 ;
         LAYER MET3 ;
         RECT  0.0 722.2 899.4 722.76 ;
         LAYER MET4 ;
         RECT  87.4 0.0 87.96 976.68 ;
         LAYER MET3 ;
         RECT  0.0 159.16 899.4 159.72 ;
         LAYER MET4 ;
         RECT  153.64 0.0 154.2 976.68 ;
         LAYER MET4 ;
         RECT  127.88 0.0 128.44 976.68 ;
         LAYER MET4 ;
         RECT  63.48 0.0 64.04 976.68 ;
         LAYER MET4 ;
         RECT  727.72 0.0 728.28 976.68 ;
         LAYER MET3 ;
         RECT  0.0 43.24 899.4 43.8 ;
         LAYER MET3 ;
         RECT  780.16 203.32 899.4 203.88 ;
         LAYER MET3 ;
         RECT  731.4 790.28 899.4 790.84 ;
         LAYER MET4 ;
         RECT  8.28 0.0 8.84 976.68 ;
         LAYER MET3 ;
         RECT  780.16 245.64 899.4 246.2 ;
         LAYER MET3 ;
         RECT  0.0 646.76 899.4 647.32 ;
         LAYER MET4 ;
         RECT  402.04 0.0 402.6 976.68 ;
         LAYER MET3 ;
         RECT  0.0 37.72 89.8 38.28 ;
         LAYER MET4 ;
         RECT  628.36 0.0 628.92 976.68 ;
         LAYER MET3 ;
         RECT  716.68 882.28 899.4 882.84 ;
         LAYER MET3 ;
         RECT  0.0 184.92 117.4 185.48 ;
         LAYER MET3 ;
         RECT  0.0 609.96 899.4 610.52 ;
         LAYER MET3 ;
         RECT  96.6 321.08 899.4 321.64 ;
         LAYER MET3 ;
         RECT  0.0 199.64 899.4 200.2 ;
         LAYER MET4 ;
         RECT  149.96 0.0 150.52 976.68 ;
         LAYER MET4 ;
         RECT  814.2 0.0 814.76 976.68 ;
         LAYER MET4 ;
         RECT  884.12 0.0 884.68 976.68 ;
         LAYER MET3 ;
         RECT  0.0 477.48 899.4 478.04 ;
         LAYER MET4 ;
         RECT  793.96 0.0 794.52 976.68 ;
         LAYER MET4 ;
         RECT  260.36 6.44 260.92 976.68 ;
         LAYER MET4 ;
         RECT  446.2 0.0 446.76 976.68 ;
         LAYER MET4 ;
         RECT  457.24 0.0 457.8 976.68 ;
         LAYER MET4 ;
         RECT  56.12 0.0 56.68 976.68 ;
         LAYER MET3 ;
         RECT  733.24 218.04 899.4 218.6 ;
         LAYER MET3 ;
         RECT  721.28 48.76 899.4 49.32 ;
         LAYER MET3 ;
         RECT  80.04 319.24 899.4 319.8 ;
         LAYER MET3 ;
         RECT  755.32 490.36 899.4 490.92 ;
         LAYER MET4 ;
         RECT  483.0 0.0 483.56 976.68 ;
         LAYER MET3 ;
         RECT  0.0 898.84 899.4 899.4 ;
         LAYER MET3 ;
         RECT  0.0 282.44 117.4 283.0 ;
         LAYER MET4 ;
         RECT  416.76 20.24 417.32 976.68 ;
         LAYER MET3 ;
         RECT  0.0 146.28 899.4 146.84 ;
         LAYER MET4 ;
         RECT  321.08 12.88 321.64 976.68 ;
         LAYER MET3 ;
         RECT  0.0 823.4 899.4 823.96 ;
         LAYER MET3 ;
         RECT  892.4 889.64 899.4 890.2 ;
         LAYER MET4 ;
         RECT  297.16 0.0 297.72 976.68 ;
         LAYER MET4 ;
         RECT  764.52 0.0 765.08 976.68 ;
         LAYER MET3 ;
         RECT  716.68 545.56 899.4 546.12 ;
         LAYER MET3 ;
         RECT  398.36 0.92 899.4 1.48 ;
         LAYER MET4 ;
         RECT  427.8 0.0 428.36 976.68 ;
         LAYER MET3 ;
         RECT  716.68 856.52 899.4 857.08 ;
         LAYER MET3 ;
         RECT  655.04 10.12 899.4 10.68 ;
         LAYER MET3 ;
         RECT  0.0 495.88 177.2 496.44 ;
         LAYER MET4 ;
         RECT  387.32 0.0 387.88 5.16 ;
         LAYER MET4 ;
         RECT  115.0 0.0 115.56 976.68 ;
         LAYER MET4 ;
         RECT  254.84 0.0 255.4 5.16 ;
         LAYER MET3 ;
         RECT  95.68 311.88 899.4 312.44 ;
         LAYER MET4 ;
         RECT  240.12 0.0 240.68 976.68 ;
         LAYER MET3 ;
         RECT  0.0 241.96 100.84 242.52 ;
         LAYER MET3 ;
         RECT  716.68 234.6 899.4 235.16 ;
         LAYER MET3 ;
         RECT  780.16 260.36 899.4 260.92 ;
         LAYER MET4 ;
         RECT  113.16 0.0 113.72 976.68 ;
         LAYER MET4 ;
         RECT  286.12 0.0 286.68 976.68 ;
         LAYER MET4 ;
         RECT  595.24 0.0 595.8 976.68 ;
         LAYER MET4 ;
         RECT  424.12 0.0 424.68 976.68 ;
         LAYER MET4 ;
         RECT  563.96 0.0 564.52 976.68 ;
         LAYER MET4 ;
         RECT  370.76 0.0 371.32 5.16 ;
         LAYER MET3 ;
         RECT  0.0 402.04 899.4 402.6 ;
         LAYER MET3 ;
         RECT  0.0 240.12 160.64 240.68 ;
         LAYER MET4 ;
         RECT  836.28 0.0 836.84 976.68 ;
         LAYER MET4 ;
         RECT  839.96 0.0 840.52 976.68 ;
         LAYER MET4 ;
         RECT  324.76 0.0 325.32 976.68 ;
         LAYER MET3 ;
         RECT  0.0 238.28 899.4 238.84 ;
         LAYER MET4 ;
         RECT  337.64 0.0 338.2 5.16 ;
         LAYER MET4 ;
         RECT  120.52 0.0 121.08 976.68 ;
         LAYER MET4 ;
         RECT  85.56 0.0 86.12 976.68 ;
         LAYER MET4 ;
         RECT  545.56 0.0 546.12 976.68 ;
         LAYER MET4 ;
         RECT  218.04 0.0 218.6 976.68 ;
         LAYER MET4 ;
         RECT  508.76 0.0 509.32 976.68 ;
         LAYER MET3 ;
         RECT  0.0 576.84 899.4 577.4 ;
         LAYER MET3 ;
         RECT  0.0 847.32 899.4 847.88 ;
         LAYER MET4 ;
         RECT  175.72 0.0 176.28 976.68 ;
         LAYER MET3 ;
         RECT  716.68 633.88 899.4 634.44 ;
         LAYER MET3 ;
         RECT  655.04 11.96 899.4 12.52 ;
         LAYER MET3 ;
         RECT  0.0 974.28 899.4 974.84 ;
         LAYER MET4 ;
         RECT  874.92 0.0 875.48 976.68 ;
         LAYER MET3 ;
         RECT  0.0 817.88 899.4 818.44 ;
         LAYER MET3 ;
         RECT  0.0 965.08 899.4 965.64 ;
         LAYER MET3 ;
         RECT  687.24 28.52 899.4 29.08 ;
         LAYER MET3 ;
         RECT  0.0 120.52 117.4 121.08 ;
         LAYER MET4 ;
         RECT  221.72 12.88 222.28 976.68 ;
         LAYER MET4 ;
         RECT  238.28 14.72 238.84 976.68 ;
         LAYER MET3 ;
         RECT  755.32 639.4 899.4 639.96 ;
         LAYER MET4 ;
         RECT  370.76 18.4 371.32 976.68 ;
         LAYER MET4 ;
         RECT  503.24 0.0 503.8 976.68 ;
         LAYER MET3 ;
         RECT  0.0 379.96 899.4 380.52 ;
         LAYER MET3 ;
         RECT  780.16 179.4 899.4 179.96 ;
         LAYER MET3 ;
         RECT  0.0 92.92 100.84 93.48 ;
         LAYER MET4 ;
         RECT  703.8 0.0 704.36 976.68 ;
         LAYER MET4 ;
         RECT  827.08 0.0 827.64 976.68 ;
         LAYER MET3 ;
         RECT  810.52 946.68 899.4 947.24 ;
         LAYER MET4 ;
         RECT  444.36 0.0 444.92 976.68 ;
         LAYER MET4 ;
         RECT  806.84 0.0 807.4 976.68 ;
         LAYER MET3 ;
         RECT  0.0 6.44 110.04 7.0 ;
         LAYER MET3 ;
         RECT  0.0 529.0 899.4 529.56 ;
         LAYER MET3 ;
         RECT  38.64 50.6 899.4 51.16 ;
         LAYER MET4 ;
         RECT  385.48 0.0 386.04 976.68 ;
         LAYER MET3 ;
         RECT  780.16 96.6 899.4 97.16 ;
         LAYER MET3 ;
         RECT  0.0 503.24 899.4 503.8 ;
         LAYER MET3 ;
         RECT  0.0 836.28 899.4 836.84 ;
         LAYER MET3 ;
         RECT  0.0 788.44 142.24 789.0 ;
         LAYER MET3 ;
         RECT  0.0 856.52 177.2 857.08 ;
         LAYER MET4 ;
         RECT  632.04 0.0 632.6 976.68 ;
         LAYER MET3 ;
         RECT  0.0 162.84 899.4 163.4 ;
         LAYER MET3 ;
         RECT  132.48 23.0 899.4 23.56 ;
         LAYER MET4 ;
         RECT  709.32 0.0 709.88 976.68 ;
         LAYER MET3 ;
         RECT  93.84 295.32 899.4 295.88 ;
         LAYER MET3 ;
         RECT  0.0 558.44 177.2 559.0 ;
         LAYER MET4 ;
         RECT  230.92 0.0 231.48 976.68 ;
         LAYER MET4 ;
         RECT  254.84 12.88 255.4 976.68 ;
         LAYER MET3 ;
         RECT  0.0 245.64 117.4 246.2 ;
         LAYER MET3 ;
         RECT  132.48 39.56 899.4 40.12 ;
         LAYER MET3 ;
         RECT  0.0 790.28 162.48 790.84 ;
         LAYER MET4 ;
         RECT  687.24 20.24 687.8 976.68 ;
         LAYER MET3 ;
         RECT  92.92 293.48 899.4 294.04 ;
         LAYER MET4 ;
         RECT  828.92 0.0 829.48 976.68 ;
         LAYER MET3 ;
         RECT  716.68 670.68 899.4 671.24 ;
         LAYER MET4 ;
         RECT  738.76 0.0 739.32 976.68 ;
         LAYER MET4 ;
         RECT  186.76 0.0 187.32 976.68 ;
         LAYER MET4 ;
         RECT  188.6 0.0 189.16 5.16 ;
         LAYER MET3 ;
         RECT  0.0 944.84 899.4 945.4 ;
         LAYER MET4 ;
         RECT  0.92 0.0 1.48 54.84 ;
         LAYER MET4 ;
         RECT  803.16 0.0 803.72 976.68 ;
         LAYER MET4 ;
         RECT  729.56 0.0 730.12 976.68 ;
         LAYER MET3 ;
         RECT  716.68 657.8 899.4 658.36 ;
         LAYER MET4 ;
         RECT  343.16 6.44 343.72 976.68 ;
         LAYER MET3 ;
         RECT  0.0 749.8 899.4 750.36 ;
         LAYER MET3 ;
         RECT  0.0 755.32 899.4 755.88 ;
         LAYER MET4 ;
         RECT  484.84 0.0 485.4 15.28 ;
         LAYER MET4 ;
         RECT  790.28 0.0 790.84 976.68 ;
         LAYER MET3 ;
         RECT  0.0 887.8 142.24 888.36 ;
         LAYER MET4 ;
         RECT  350.52 0.0 351.08 976.68 ;
         LAYER MET4 ;
         RECT  713.0 0.0 713.56 976.68 ;
         LAYER MET4 ;
         RECT  624.68 0.0 625.24 976.68 ;
         LAYER MET4 ;
         RECT  825.24 0.0 825.8 976.68 ;
         LAYER MET4 ;
         RECT  843.64 0.0 844.2 976.68 ;
         LAYER MET3 ;
         RECT  0.0 157.32 899.4 157.88 ;
         LAYER MET4 ;
         RECT  103.96 0.0 104.52 976.68 ;
         LAYER MET3 ;
         RECT  0.0 149.96 899.4 150.52 ;
         LAYER MET3 ;
         RECT  0.0 659.64 899.4 660.2 ;
         LAYER MET3 ;
         RECT  0.0 972.44 741.16 973.0 ;
         LAYER MET4 ;
         RECT  817.88 0.0 818.44 976.68 ;
         LAYER MET3 ;
         RECT  0.0 565.8 160.64 566.36 ;
         LAYER MET3 ;
         RECT  780.16 282.44 899.4 283.0 ;
         LAYER MET4 ;
         RECT  23.0 0.0 23.56 976.68 ;
         LAYER MET3 ;
         RECT  870.32 954.04 899.4 954.6 ;
         LAYER MET3 ;
         RECT  0.0 471.96 177.2 472.52 ;
         LAYER MET4 ;
         RECT  48.76 0.0 49.32 976.68 ;
         LAYER MET3 ;
         RECT  0.0 514.28 142.24 514.84 ;
         LAYER MET4 ;
         RECT  135.24 0.0 135.8 976.68 ;
         LAYER MET4 ;
         RECT  376.28 0.0 376.84 976.68 ;
         LAYER MET4 ;
         RECT  304.52 16.56 305.08 976.68 ;
         LAYER MET4 ;
         RECT  551.08 0.0 551.64 15.28 ;
         LAYER MET4 ;
         RECT  880.44 0.0 881.0 976.68 ;
         LAYER MET3 ;
         RECT  586.96 13.8 899.4 14.36 ;
         LAYER MET4 ;
         RECT  10.12 0.0 10.68 976.68 ;
         LAYER MET3 ;
         RECT  0.0 446.2 177.2 446.76 ;
         LAYER MET3 ;
         RECT  0.0 865.72 899.4 866.28 ;
         LAYER MET4 ;
         RECT  644.92 0.0 645.48 976.68 ;
         LAYER MET4 ;
         RECT  188.6 12.88 189.16 976.68 ;
         LAYER MET3 ;
         RECT  0.0 74.52 899.4 75.08 ;
         LAYER MET3 ;
         RECT  0.0 922.76 882.84 923.32 ;
         LAYER MET4 ;
         RECT  540.04 0.0 540.6 976.68 ;
         LAYER MET3 ;
         RECT  0.0 604.44 899.4 605.0 ;
         LAYER MET4 ;
         RECT  762.68 0.0 763.24 976.68 ;
         LAYER MET4 ;
         RECT  372.6 0.0 373.16 976.68 ;
         LAYER MET4 ;
         RECT  698.28 0.0 698.84 976.68 ;
         LAYER MET4 ;
         RECT  747.96 0.0 748.52 976.68 ;
         LAYER MET3 ;
         RECT  780.16 197.8 899.4 198.36 ;
         LAYER MET3 ;
         RECT  0.0 490.36 142.24 490.92 ;
         LAYER MET4 ;
         RECT  654.12 20.24 654.68 976.68 ;
         LAYER MET4 ;
         RECT  849.16 0.0 849.72 976.68 ;
         LAYER MET4 ;
         RECT  613.64 0.0 614.2 976.68 ;
         LAYER MET4 ;
         RECT  190.44 0.0 191.0 976.68 ;
         LAYER MET4 ;
         RECT  321.08 0.0 321.64 5.16 ;
         LAYER MET4 ;
         RECT  580.52 0.0 581.08 976.68 ;
         LAYER MET3 ;
         RECT  0.0 779.24 899.4 779.8 ;
         LAYER MET4 ;
         RECT  335.8 0.0 336.36 976.68 ;
         LAYER MET3 ;
         RECT  0.0 195.96 117.4 196.52 ;
         LAYER MET4 ;
         RECT  70.84 0.0 71.4 976.68 ;
         LAYER MET4 ;
         RECT  488.52 0.0 489.08 976.68 ;
         LAYER MET4 ;
         RECT  856.52 0.0 857.08 976.68 ;
         LAYER MET3 ;
         RECT  0.0 724.04 899.4 724.6 ;
         LAYER MET3 ;
         RECT  0.0 413.08 899.4 413.64 ;
         LAYER MET3 ;
         RECT  0.0 13.8 22.64 14.36 ;
         LAYER MET4 ;
         RECT  665.16 0.0 665.72 976.68 ;
         LAYER MET3 ;
         RECT  0.0 172.04 117.4 172.6 ;
         LAYER MET3 ;
         RECT  0.0 505.08 899.4 505.64 ;
         LAYER MET4 ;
         RECT  365.24 0.0 365.8 976.68 ;
         LAYER MET3 ;
         RECT  0.0 39.56 121.08 40.12 ;
         LAYER MET4 ;
         RECT  249.32 0.0 249.88 976.68 ;
         LAYER MET4 ;
         RECT  860.2 0.0 860.76 976.68 ;
         LAYER MET4 ;
         RECT  873.08 0.0 873.64 976.68 ;
         LAYER MET3 ;
         RECT  0.0 549.24 899.4 549.8 ;
         LAYER MET4 ;
         RECT  676.2 0.0 676.76 976.68 ;
         LAYER MET4 ;
         RECT  273.24 0.0 273.8 976.68 ;
         LAYER MET4 ;
         RECT  648.6 0.0 649.16 976.68 ;
         LAYER MET3 ;
         RECT  0.0 326.6 899.4 327.16 ;
         LAYER MET3 ;
         RECT  780.16 269.56 899.4 270.12 ;
         LAYER MET3 ;
         RECT  780.16 135.24 899.4 135.8 ;
         LAYER MET3 ;
         RECT  0.0 462.76 899.4 463.32 ;
         LAYER MET4 ;
         RECT  207.0 0.0 207.56 976.68 ;
         LAYER MET4 ;
         RECT  755.32 0.0 755.88 976.68 ;
         LAYER MET3 ;
         RECT  0.0 424.12 899.4 424.68 ;
         LAYER MET3 ;
         RECT  0.0 357.88 899.4 358.44 ;
         LAYER MET3 ;
         RECT  0.0 72.68 158.8 73.24 ;
         LAYER MET3 ;
         RECT  780.16 129.72 899.4 130.28 ;
         LAYER MET3 ;
         RECT  0.0 26.68 899.4 27.24 ;
         LAYER MET3 ;
         RECT  755.32 613.64 899.4 614.2 ;
         LAYER MET4 ;
         RECT  330.28 0.0 330.84 976.68 ;
         LAYER MET4 ;
         RECT  582.36 0.0 582.92 976.68 ;
         LAYER MET3 ;
         RECT  0.0 317.4 160.64 317.96 ;
         LAYER MET3 ;
         RECT  755.32 689.08 899.4 689.64 ;
         LAYER MET4 ;
         RECT  525.32 0.0 525.88 976.68 ;
         LAYER MET3 ;
         RECT  716.68 558.44 899.4 559.0 ;
         LAYER MET4 ;
         RECT  470.12 0.0 470.68 976.68 ;
         LAYER MET3 ;
         RECT  892.4 906.2 899.4 906.76 ;
         LAYER MET3 ;
         RECT  0.0 251.16 899.4 251.72 ;
         LAYER MET4 ;
         RECT  131.56 0.0 132.12 976.68 ;
         LAYER MET3 ;
         RECT  780.16 207.0 899.4 207.56 ;
         LAYER MET3 ;
         RECT  0.0 600.76 899.4 601.32 ;
         LAYER MET3 ;
         RECT  0.0 50.6 7.0 51.16 ;
         LAYER MET3 ;
         RECT  0.0 385.48 899.4 386.04 ;
         LAYER MET4 ;
         RECT  779.24 0.0 779.8 976.68 ;
         LAYER MET3 ;
         RECT  0.0 161.0 177.2 161.56 ;
         LAYER MET3 ;
         RECT  716.68 322.92 899.4 323.48 ;
         LAYER MET3 ;
         RECT  80.04 302.68 899.4 303.24 ;
         LAYER MET3 ;
         RECT  0.0 422.28 177.2 422.84 ;
         LAYER MET3 ;
         RECT  0.0 714.84 142.24 715.4 ;
         LAYER MET3 ;
         RECT  780.16 195.96 899.4 196.52 ;
         LAYER MET4 ;
         RECT  845.48 0.0 846.04 976.68 ;
         LAYER MET3 ;
         RECT  716.68 595.24 899.4 595.8 ;
         LAYER MET3 ;
         RECT  0.0 153.64 899.4 154.2 ;
         LAYER MET4 ;
         RECT  655.96 0.0 656.52 976.68 ;
         LAYER MET3 ;
         RECT  716.68 521.64 899.4 522.2 ;
         LAYER MET4 ;
         RECT  429.64 0.0 430.2 976.68 ;
         LAYER MET4 ;
         RECT  459.08 0.0 459.64 976.68 ;
         LAYER MET4 ;
         RECT  490.36 0.0 490.92 976.68 ;
         LAYER MET3 ;
         RECT  0.0 915.4 899.4 915.96 ;
         LAYER MET4 ;
         RECT  621.0 0.0 621.56 976.68 ;
         LAYER MET3 ;
         RECT  0.0 551.08 899.4 551.64 ;
         LAYER MET3 ;
         RECT  0.0 52.44 899.4 53.0 ;
         LAYER MET4 ;
         RECT  310.04 0.0 310.6 976.68 ;
         LAYER MET3 ;
         RECT  0.0 506.92 899.4 507.48 ;
         LAYER MET3 ;
         RECT  91.08 8.28 899.4 8.84 ;
         LAYER MET3 ;
         RECT  0.0 383.64 177.2 384.2 ;
         LAYER MET3 ;
         RECT  689.08 19.32 899.4 19.88 ;
         LAYER MET3 ;
         RECT  0.0 243.8 117.4 244.36 ;
         LAYER MET4 ;
         RECT  637.56 0.0 638.12 976.68 ;
         LAYER MET3 ;
         RECT  0.0 652.28 899.4 652.84 ;
         LAYER MET3 ;
         RECT  797.64 265.88 899.4 266.44 ;
         LAYER MET3 ;
         RECT  0.0 657.8 177.2 658.36 ;
         LAYER MET3 ;
         RECT  716.68 409.4 899.4 409.96 ;
         LAYER MET3 ;
         RECT  0.0 234.6 177.2 235.16 ;
         LAYER MET4 ;
         RECT  597.08 0.0 597.64 976.68 ;
         LAYER MET4 ;
         RECT  111.32 0.0 111.88 976.68 ;
         LAYER MET4 ;
         RECT  696.44 0.0 697.0 976.68 ;
         LAYER MET3 ;
         RECT  0.0 273.24 117.4 273.8 ;
         LAYER MET3 ;
         RECT  755.32 589.72 899.4 590.28 ;
         LAYER MET4 ;
         RECT  287.96 0.0 288.52 5.16 ;
         LAYER MET3 ;
         RECT  0.0 486.68 899.4 487.24 ;
         LAYER MET3 ;
         RECT  0.0 473.8 899.4 474.36 ;
         LAYER MET4 ;
         RECT  773.72 0.0 774.28 976.68 ;
         LAYER MET4 ;
         RECT  440.68 0.0 441.24 976.68 ;
         LAYER MET3 ;
         RECT  731.4 438.84 899.4 439.4 ;
         LAYER MET4 ;
         RECT  319.24 0.0 319.8 976.68 ;
         LAYER MET3 ;
         RECT  0.0 803.16 899.4 803.72 ;
         LAYER MET3 ;
         RECT  780.16 256.68 899.4 257.24 ;
         LAYER MET4 ;
         RECT  179.4 0.0 179.96 9.76 ;
         LAYER MET4 ;
         RECT  155.48 12.88 156.04 976.68 ;
         LAYER MET4 ;
         RECT  308.2 0.0 308.76 976.68 ;
         LAYER MET3 ;
         RECT  0.0 801.32 899.4 801.88 ;
         LAYER MET4 ;
         RECT  293.48 6.44 294.04 976.68 ;
         LAYER MET4 ;
         RECT  208.84 0.0 209.4 976.68 ;
         LAYER MET4 ;
         RECT  405.72 0.0 406.28 976.68 ;
         LAYER MET3 ;
         RECT  0.0 256.68 117.4 257.24 ;
         LAYER MET3 ;
         RECT  0.0 232.76 899.4 233.32 ;
         LAYER MET3 ;
         RECT  780.16 111.32 899.4 111.88 ;
         LAYER MET3 ;
         RECT  0.0 0.92 113.72 1.48 ;
         LAYER MET3 ;
         RECT  780.16 208.84 899.4 209.4 ;
         LAYER MET3 ;
         RECT  0.0 83.72 7.0 84.28 ;
         LAYER MET3 ;
         RECT  0.0 709.32 899.4 709.88 ;
         LAYER MET3 ;
         RECT  0.0 622.84 899.4 623.4 ;
         LAYER MET3 ;
         RECT  0.0 731.4 899.4 731.96 ;
         LAYER MET3 ;
         RECT  0.0 705.64 899.4 706.2 ;
         LAYER MET3 ;
         RECT  0.0 626.52 899.4 627.08 ;
         LAYER MET4 ;
         RECT  164.68 0.0 165.24 976.68 ;
         LAYER MET3 ;
         RECT  0.0 562.12 899.4 562.68 ;
         LAYER MET4 ;
         RECT  205.16 0.0 205.72 5.16 ;
         LAYER MET3 ;
         RECT  0.0 608.12 177.2 608.68 ;
         LAYER MET3 ;
         RECT  0.0 795.8 899.4 796.36 ;
         LAYER MET4 ;
         RECT  775.56 0.0 776.12 976.68 ;
         LAYER MET3 ;
         RECT  0.0 812.36 160.64 812.92 ;
         LAYER MET3 ;
         RECT  0.0 902.52 881.0 903.08 ;
         LAYER MET4 ;
         RECT  173.88 0.0 174.44 976.68 ;
         LAYER MET4 ;
         RECT  282.44 0.0 283.0 976.68 ;
         LAYER MET3 ;
         RECT  0.0 374.44 899.4 375.0 ;
         LAYER MET3 ;
         RECT  0.0 41.4 87.96 41.96 ;
         LAYER MET4 ;
         RECT  299.0 0.0 299.56 976.68 ;
         LAYER MET4 ;
         RECT  172.04 12.88 172.6 976.68 ;
         LAYER MET3 ;
         RECT  809.6 917.24 899.4 917.8 ;
         LAYER MET3 ;
         RECT  0.0 286.12 117.4 286.68 ;
         LAYER MET4 ;
         RECT  724.04 0.0 724.6 976.68 ;
         LAYER MET3 ;
         RECT  0.0 773.72 899.4 774.28 ;
         LAYER MET3 ;
         RECT  755.32 563.96 899.4 564.52 ;
         LAYER MET3 ;
         RECT  0.0 205.16 117.4 205.72 ;
         LAYER MET4 ;
         RECT  383.64 0.0 384.2 976.68 ;
         LAYER MET4 ;
         RECT  622.84 0.0 623.4 976.68 ;
         LAYER MET3 ;
         RECT  733.24 466.44 899.4 467.0 ;
         LAYER MET3 ;
         RECT  0.0 324.76 80.6 325.32 ;
         LAYER MET4 ;
         RECT  74.52 0.0 75.08 976.68 ;
         LAYER MET3 ;
         RECT  780.16 280.6 899.4 281.16 ;
         LAYER MET3 ;
         RECT  0.0 466.44 160.64 467.0 ;
         LAYER MET3 ;
         RECT  0.0 943.0 766.0 943.56 ;
         LAYER MET3 ;
         RECT  716.68 161.0 899.4 161.56 ;
         LAYER MET3 ;
         RECT  716.68 845.48 899.4 846.04 ;
         LAYER MET4 ;
         RECT  609.96 0.0 610.52 976.68 ;
         LAYER MET4 ;
         RECT  81.88 0.0 82.44 976.68 ;
         LAYER MET3 ;
         RECT  0.0 683.56 177.2 684.12 ;
         LAYER MET3 ;
         RECT  0.0 584.2 899.4 584.76 ;
         LAYER MET4 ;
         RECT  733.24 0.0 733.8 976.68 ;
         LAYER MET3 ;
         RECT  797.64 142.6 899.4 143.16 ;
         LAYER MET3 ;
         RECT  797.64 241.96 899.4 242.52 ;
         LAYER MET3 ;
         RECT  0.0 287.96 899.4 288.52 ;
         LAYER MET3 ;
         RECT  716.68 459.08 899.4 459.64 ;
         LAYER MET3 ;
         RECT  0.0 889.64 160.64 890.2 ;
         LAYER MET3 ;
         RECT  739.68 67.16 899.4 67.72 ;
         LAYER MET4 ;
         RECT  52.44 0.0 53.0 976.68 ;
         LAYER MET4 ;
         RECT  280.6 20.24 281.16 976.68 ;
         LAYER MET3 ;
         RECT  0.0 876.76 881.0 877.32 ;
         LAYER MET4 ;
         RECT  736.92 0.0 737.48 976.68 ;
         LAYER MET3 ;
         RECT  0.0 264.04 899.4 264.6 ;
         LAYER MET3 ;
         RECT  0.0 882.28 177.2 882.84 ;
         LAYER MET4 ;
         RECT  201.48 0.0 202.04 976.68 ;
         LAYER MET4 ;
         RECT  192.28 0.0 192.84 976.68 ;
         LAYER MET3 ;
         RECT  0.0 214.36 899.4 214.92 ;
         LAYER MET3 ;
         RECT  739.68 72.68 899.4 73.24 ;
         LAYER MET3 ;
         RECT  0.0 425.96 899.4 426.52 ;
         LAYER MET4 ;
         RECT  172.04 0.0 172.6 5.16 ;
         LAYER MET4 ;
         RECT  562.12 0.0 562.68 976.68 ;
         LAYER MET4 ;
         RECT  32.2 0.0 32.76 976.68 ;
         LAYER MET3 ;
         RECT  0.0 508.76 177.2 509.32 ;
         LAYER MET4 ;
         RECT  788.44 0.0 789.0 976.68 ;
         LAYER MET3 ;
         RECT  0.0 308.2 80.6 308.76 ;
         LAYER MET3 ;
         RECT  0.0 455.4 899.4 455.96 ;
         LAYER MET3 ;
         RECT  0.0 32.2 899.4 32.76 ;
         LAYER MET3 ;
         RECT  821.56 46.92 899.4 47.48 ;
         LAYER MET3 ;
         RECT  19.32 113.16 899.4 113.72 ;
         LAYER MET3 ;
         RECT  716.68 124.2 899.4 124.76 ;
         LAYER MET3 ;
         RECT  733.24 339.48 899.4 340.04 ;
         LAYER MET4 ;
         RECT  598.92 0.0 599.48 976.68 ;
         LAYER MET4 ;
         RECT  744.28 0.0 744.84 976.68 ;
         LAYER MET3 ;
         RECT  780.16 122.36 899.4 122.92 ;
         LAYER MET3 ;
         RECT  0.0 742.44 899.4 743.0 ;
         LAYER MET3 ;
         RECT  0.0 746.12 899.4 746.68 ;
         LAYER MET3 ;
         RECT  0.0 21.16 32.76 21.72 ;
         LAYER MET4 ;
         RECT  326.6 0.0 327.16 976.68 ;
         LAYER MET4 ;
         RECT  414.92 0.0 415.48 976.68 ;
         LAYER MET4 ;
         RECT  670.68 0.0 671.24 976.68 ;
         LAYER MET3 ;
         RECT  0.0 137.08 899.4 137.64 ;
         LAYER MET3 ;
         RECT  0.0 545.56 177.2 546.12 ;
         LAYER MET3 ;
         RECT  0.0 707.48 177.2 708.04 ;
         LAYER MET4 ;
         RECT  477.48 0.0 478.04 976.68 ;
         LAYER MET3 ;
         RECT  716.68 422.28 899.4 422.84 ;
         LAYER MET4 ;
         RECT  869.4 0.0 869.96 976.68 ;
         LAYER MET4 ;
         RECT  468.28 0.0 468.84 976.68 ;
         LAYER MET3 ;
         RECT  716.68 733.24 899.4 733.8 ;
         LAYER MET3 ;
         RECT  0.0 183.08 117.4 183.64 ;
         LAYER MET4 ;
         RECT  354.2 0.0 354.76 5.16 ;
         LAYER MET4 ;
         RECT  407.56 0.0 408.12 976.68 ;
         LAYER MET4 ;
         RECT  600.76 0.0 601.32 976.68 ;
         LAYER MET3 ;
         RECT  0.0 926.44 740.24 927.0 ;
         LAYER MET4 ;
         RECT  345.0 0.0 345.56 976.68 ;
         LAYER MET4 ;
         RECT  328.44 0.0 329.0 976.68 ;
         LAYER MET3 ;
         RECT  755.32 440.68 899.4 441.24 ;
         LAYER MET3 ;
         RECT  0.0 354.2 899.4 354.76 ;
         LAYER MET3 ;
         RECT  80.04 330.28 899.4 330.84 ;
         LAYER MET4 ;
         RECT  630.2 0.0 630.76 976.68 ;
         LAYER MET3 ;
         RECT  0.0 858.36 899.4 858.92 ;
         LAYER MET4 ;
         RECT  760.84 0.0 761.4 976.68 ;
         LAYER MET3 ;
         RECT  0.0 218.04 160.64 218.6 ;
         LAYER MET3 ;
         RECT  0.0 573.16 899.4 573.72 ;
         LAYER MET4 ;
         RECT  129.72 0.0 130.28 976.68 ;
         LAYER MET4 ;
         RECT  245.64 0.0 246.2 962.88 ;
         LAYER MET4 ;
         RECT  359.72 6.44 360.28 976.68 ;
         LAYER MET4 ;
         RECT  876.76 0.0 877.32 976.68 ;
         LAYER MET3 ;
         RECT  0.0 15.64 271.04 16.2 ;
         LAYER MET3 ;
         RECT  0.0 361.56 899.4 362.12 ;
         LAYER MET4 ;
         RECT  223.56 0.0 224.12 976.68 ;
         LAYER MET3 ;
         RECT  0.0 115.0 899.4 115.56 ;
         LAYER MET3 ;
         RECT  0.0 602.6 899.4 603.16 ;
         LAYER MET3 ;
         RECT  0.0 453.56 899.4 454.12 ;
         LAYER MET4 ;
         RECT  786.6 0.0 787.16 976.68 ;
         LAYER MET4 ;
         RECT  832.6 0.0 833.16 976.68 ;
         LAYER MET3 ;
         RECT  797.64 116.84 899.4 117.4 ;
         LAYER MET3 ;
         RECT  0.0 299.0 899.4 299.56 ;
         LAYER MET3 ;
         RECT  0.0 94.76 117.4 95.32 ;
         LAYER MET4 ;
         RECT  197.8 0.0 198.36 976.68 ;
         LAYER MET3 ;
         RECT  0.0 229.08 899.4 229.64 ;
         LAYER MET3 ;
         RECT  733.24 812.36 899.4 812.92 ;
         LAYER MET3 ;
         RECT  0.0 170.2 117.4 170.76 ;
         LAYER MET3 ;
         RECT  0.0 678.04 899.4 678.6 ;
         LAYER MET3 ;
         RECT  0.0 878.6 899.4 879.16 ;
         LAYER MET3 ;
         RECT  0.0 460.92 899.4 461.48 ;
         LAYER MET3 ;
         RECT  0.0 126.04 899.4 126.6 ;
         LAYER MET3 ;
         RECT  0.0 571.32 177.2 571.88 ;
         LAYER MET3 ;
         RECT  0.0 124.2 177.2 124.76 ;
         LAYER MET3 ;
         RECT  0.0 643.08 899.4 643.64 ;
         LAYER MET3 ;
         RECT  810.52 930.12 899.4 930.68 ;
         LAYER MET4 ;
         RECT  547.4 0.0 547.96 976.68 ;
         LAYER MET3 ;
         RECT  0.0 155.48 899.4 156.04 ;
         LAYER MET4 ;
         RECT  26.68 0.0 27.24 976.68 ;
         LAYER MET3 ;
         RECT  0.0 589.72 142.24 590.28 ;
         LAYER MET3 ;
         RECT  716.68 869.4 899.4 869.96 ;
         LAYER MET4 ;
         RECT  586.04 20.24 586.6 976.68 ;
         LAYER MET3 ;
         RECT  716.68 495.88 899.4 496.44 ;
         LAYER MET3 ;
         RECT  0.0 845.48 177.2 846.04 ;
         LAYER MET3 ;
         RECT  0.0 168.36 117.4 168.92 ;
         LAYER MET4 ;
         RECT  43.24 0.0 43.8 976.68 ;
         LAYER MET3 ;
         RECT  0.0 799.48 899.4 800.04 ;
         LAYER MET3 ;
         RECT  0.0 433.32 899.4 433.88 ;
         LAYER MET3 ;
         RECT  716.68 720.36 899.4 720.92 ;
         LAYER MET4 ;
         RECT  333.96 0.0 334.52 976.68 ;
         LAYER MET3 ;
         RECT  817.88 41.4 899.4 41.96 ;
         LAYER MET3 ;
         RECT  0.0 884.12 881.0 884.68 ;
         LAYER MET3 ;
         RECT  0.0 698.28 899.4 698.84 ;
         LAYER MET4 ;
         RECT  751.64 0.0 752.2 976.68 ;
         LAYER MET4 ;
         RECT  556.6 0.0 557.16 976.68 ;
         LAYER MET4 ;
         RECT  770.04 0.0 770.6 970.24 ;
         LAYER MET3 ;
         RECT  0.0 895.16 177.2 895.72 ;
         LAYER MET4 ;
         RECT  858.36 0.0 858.92 976.68 ;
         LAYER MET3 ;
         RECT  780.16 181.24 899.4 181.8 ;
         LAYER MET4 ;
         RECT  118.68 0.0 119.24 976.68 ;
         LAYER MET3 ;
         RECT  0.0 431.48 899.4 432.04 ;
         LAYER MET3 ;
         RECT  0.0 300.84 899.4 301.4 ;
         LAYER MET4 ;
         RECT  433.32 0.0 433.88 976.68 ;
         LAYER MET4 ;
         RECT  148.12 0.0 148.68 976.68 ;
         LAYER MET3 ;
         RECT  0.0 140.76 160.64 141.32 ;
         LAYER MET4 ;
         RECT  194.12 6.44 194.68 976.68 ;
         LAYER MET3 ;
         RECT  716.68 683.56 899.4 684.12 ;
         LAYER MET3 ;
         RECT  0.0 692.76 899.4 693.32 ;
         LAYER MET3 ;
         RECT  733.24 367.08 899.4 367.64 ;
         LAYER MET3 ;
         RECT  0.0 700.12 899.4 700.68 ;
         LAYER MET4 ;
         RECT  400.2 0.0 400.76 976.68 ;
         LAYER MET4 ;
         RECT  674.36 0.0 674.92 976.68 ;
         LAYER MET4 ;
         RECT  253.0 0.0 253.56 976.68 ;
         LAYER MET3 ;
         RECT  716.68 223.56 899.4 224.12 ;
         LAYER MET3 ;
         RECT  733.24 140.76 899.4 141.32 ;
         LAYER MET3 ;
         RECT  0.0 254.84 117.4 255.4 ;
         LAYER MET3 ;
         RECT  0.0 201.48 899.4 202.04 ;
         LAYER MET3 ;
         RECT  817.88 76.36 899.4 76.92 ;
         LAYER MET3 ;
         RECT  0.0 479.32 899.4 479.88 ;
         LAYER MET4 ;
         RECT  140.76 0.0 141.32 976.68 ;
         LAYER MET3 ;
         RECT  0.0 346.84 177.2 347.4 ;
         LAYER MET4 ;
         RECT  494.04 0.0 494.6 976.68 ;
         LAYER MET4 ;
         RECT  690.92 0.0 691.48 976.68 ;
         LAYER MET4 ;
         RECT  841.8 0.0 842.36 976.68 ;
         LAYER MET4 ;
         RECT  24.84 0.0 25.4 976.68 ;
         LAYER MET4 ;
         RECT  558.44 0.0 559.0 976.68 ;
         LAYER MET4 ;
         RECT  471.96 0.0 472.52 976.68 ;
         LAYER MET4 ;
         RECT  363.4 0.0 363.96 976.68 ;
         LAYER MET4 ;
         RECT  523.48 0.0 524.04 976.68 ;
         LAYER MET3 ;
         RECT  780.16 131.56 899.4 132.12 ;
         LAYER MET3 ;
         RECT  0.0 764.52 142.24 765.08 ;
         LAYER MET3 ;
         RECT  755.32 414.92 899.4 415.48 ;
         LAYER MET3 ;
         RECT  755.32 764.52 899.4 765.08 ;
         LAYER MET4 ;
         RECT  352.36 0.0 352.92 976.68 ;
         LAYER MET4 ;
         RECT  170.2 0.0 170.76 976.68 ;
         LAYER MET3 ;
         RECT  733.24 713.0 899.4 713.56 ;
         LAYER MET3 ;
         RECT  0.0 805.0 899.4 805.56 ;
         LAYER MET4 ;
         RECT  30.36 0.0 30.92 976.68 ;
         LAYER MET3 ;
         RECT  0.0 641.24 899.4 641.8 ;
         LAYER MET3 ;
         RECT  866.64 950.36 899.4 950.92 ;
         LAYER MET4 ;
         RECT  124.2 0.0 124.76 976.68 ;
         LAYER MET3 ;
         RECT  552.92 15.64 899.4 16.2 ;
         LAYER MET4 ;
         RECT  157.32 0.0 157.88 976.68 ;
         LAYER MET3 ;
         RECT  0.0 871.24 882.84 871.8 ;
         LAYER MET3 ;
         RECT  0.0 216.2 100.84 216.76 ;
         LAYER MET3 ;
         RECT  0.0 701.96 899.4 702.52 ;
         LAYER MET3 ;
         RECT  0.0 133.4 117.4 133.96 ;
         LAYER MET3 ;
         RECT  780.16 98.44 899.4 99.0 ;
         LAYER MET3 ;
         RECT  0.0 632.04 899.4 632.6 ;
         LAYER MET3 ;
         RECT  0.0 873.08 899.4 873.64 ;
         LAYER MET4 ;
         RECT  391.0 0.0 391.56 976.68 ;
         LAYER MET4 ;
         RECT  13.8 0.0 14.36 976.68 ;
         LAYER MET3 ;
         RECT  869.4 943.0 899.4 943.56 ;
         LAYER MET3 ;
         RECT  0.0 552.92 899.4 553.48 ;
         LAYER MET3 ;
         RECT  733.24 91.08 899.4 91.64 ;
         LAYER MET3 ;
         RECT  0.0 175.72 899.4 176.28 ;
         LAYER MET3 ;
         RECT  780.16 103.96 899.4 104.52 ;
         LAYER MET3 ;
         RECT  0.0 109.48 117.4 110.04 ;
         LAYER MET3 ;
         RECT  780.16 258.52 899.4 259.08 ;
         LAYER MET3 ;
         RECT  0.0 753.48 899.4 754.04 ;
         LAYER MET4 ;
         RECT  821.56 71.76 822.12 976.68 ;
         LAYER MET3 ;
         RECT  0.0 370.76 899.4 371.32 ;
         LAYER MET3 ;
         RECT  755.32 341.32 899.4 341.88 ;
         LAYER MET3 ;
         RECT  0.0 725.88 899.4 726.44 ;
         LAYER MET4 ;
         RECT  481.16 0.0 481.72 976.68 ;
         LAYER MET3 ;
         RECT  0.0 407.56 899.4 408.12 ;
         LAYER MET4 ;
         RECT  878.6 0.0 879.16 976.68 ;
         LAYER MET4 ;
         RECT  687.24 0.0 687.8 17.12 ;
         LAYER MET3 ;
         RECT  733.24 565.8 899.4 566.36 ;
         LAYER MET3 ;
         RECT  731.4 690.92 899.4 691.48 ;
         LAYER MET3 ;
         RECT  0.0 650.44 899.4 651.0 ;
         LAYER MET4 ;
         RECT  389.16 0.0 389.72 976.68 ;
         LAYER MET4 ;
         RECT  392.84 0.0 393.4 976.68 ;
         LAYER MET4 ;
         RECT  403.88 20.24 404.44 976.68 ;
         LAYER MET3 ;
         RECT  877.68 957.72 899.4 958.28 ;
         LAYER MET4 ;
         RECT  589.72 0.0 590.28 976.68 ;
         LAYER MET4 ;
         RECT  346.84 0.0 347.4 976.68 ;
         LAYER MET4 ;
         RECT  0.92 114.08 1.48 976.68 ;
         LAYER MET4 ;
         RECT  11.96 0.0 12.52 976.68 ;
         LAYER MET3 ;
         RECT  0.0 262.2 899.4 262.76 ;
         LAYER MET3 ;
         RECT  0.0 841.8 899.4 842.36 ;
         LAYER MET4 ;
         RECT  578.68 0.0 579.24 976.68 ;
         LAYER MET4 ;
         RECT  705.64 0.0 706.2 976.68 ;
         LAYER MET4 ;
         RECT  473.8 0.0 474.36 976.68 ;
         LAYER MET4 ;
         RECT  871.24 0.0 871.8 976.68 ;
         LAYER MET3 ;
         RECT  0.0 814.2 142.24 814.76 ;
         LAYER MET4 ;
         RECT  92.92 0.0 93.48 976.68 ;
         LAYER MET4 ;
         RECT  484.84 20.24 485.4 976.68 ;
         LAYER MET3 ;
         RECT  0.0 475.64 899.4 476.2 ;
         LAYER MET4 ;
         RECT  576.84 0.0 577.4 976.68 ;
         LAYER MET4 ;
         RECT  80.04 0.0 80.6 976.68 ;
         LAYER MET3 ;
         RECT  716.68 383.64 899.4 384.2 ;
         LAYER MET4 ;
         RECT  679.88 0.0 680.44 976.68 ;
         LAYER MET3 ;
         RECT  0.0 470.12 899.4 470.68 ;
         LAYER MET4 ;
         RECT  532.68 0.0 533.24 976.68 ;
         LAYER MET3 ;
         RECT  0.0 494.04 899.4 494.6 ;
         LAYER MET3 ;
         RECT  0.0 615.48 142.24 616.04 ;
         LAYER MET4 ;
         RECT  801.32 0.0 801.88 976.68 ;
         LAYER MET3 ;
         RECT  0.0 46.92 800.04 47.48 ;
         LAYER MET4 ;
         RECT  854.68 0.0 855.24 976.68 ;
         LAYER MET3 ;
         RECT  0.0 806.84 177.2 807.4 ;
         LAYER MET3 ;
         RECT  0.0 613.64 142.24 614.2 ;
         LAYER MET4 ;
         RECT  882.28 0.0 882.84 976.68 ;
         LAYER MET3 ;
         RECT  0.0 207.0 117.4 207.56 ;
         LAYER MET4 ;
         RECT  812.36 0.0 812.92 976.68 ;
         LAYER MET3 ;
         RECT  817.88 57.96 899.4 58.52 ;
         LAYER MET3 ;
         RECT  716.68 471.96 899.4 472.52 ;
         LAYER MET4 ;
         RECT  891.48 0.0 892.04 976.68 ;
         LAYER MET4 ;
         RECT  216.2 0.0 216.76 976.68 ;
         LAYER MET4 ;
         RECT  584.2 0.0 584.76 976.68 ;
         LAYER MET3 ;
         RECT  0.0 681.72 899.4 682.28 ;
         LAYER MET3 ;
         RECT  780.16 267.72 899.4 268.28 ;
         LAYER MET3 ;
         RECT  0.0 784.76 899.4 785.32 ;
         LAYER MET4 ;
         RECT  265.88 0.0 266.44 976.68 ;
         LAYER MET4 ;
         RECT  685.4 0.0 685.96 976.68 ;
         LAYER MET4 ;
         RECT  453.56 0.0 454.12 976.68 ;
         LAYER MET3 ;
         RECT  0.0 315.56 142.24 316.12 ;
         LAYER MET3 ;
         RECT  0.0 387.32 899.4 387.88 ;
         LAYER MET4 ;
         RECT  269.56 0.0 270.12 976.68 ;
         LAYER MET4 ;
         RECT  361.56 0.0 362.12 976.68 ;
         LAYER MET3 ;
         RECT  0.0 578.68 899.4 579.24 ;
         LAYER MET3 ;
         RECT  0.0 105.8 117.4 106.36 ;
         LAYER MET3 ;
         RECT  0.0 727.72 899.4 728.28 ;
         LAYER MET3 ;
         RECT  0.0 738.76 142.24 739.32 ;
         LAYER MET3 ;
         RECT  0.0 782.92 177.2 783.48 ;
         LAYER MET4 ;
         RECT  367.08 0.0 367.64 976.68 ;
         LAYER MET3 ;
         RECT  0.0 368.92 899.4 369.48 ;
         LAYER MET4 ;
         RECT  96.6 0.0 97.16 976.68 ;
         LAYER MET4 ;
         RECT  258.52 0.0 259.08 976.68 ;
         LAYER MET3 ;
         RECT  0.0 330.28 77.84 330.84 ;
         LAYER MET4 ;
         RECT  681.72 0.0 682.28 976.68 ;
         LAYER MET4 ;
         RECT  89.24 0.0 89.8 976.68 ;
         LAYER MET4 ;
         RECT  830.76 0.0 831.32 976.68 ;
         LAYER MET4 ;
         RECT  486.68 0.0 487.24 976.68 ;
         LAYER MET3 ;
         RECT  689.08 17.48 899.4 18.04 ;
         LAYER MET3 ;
         RECT  0.0 30.36 899.4 30.92 ;
         LAYER MET3 ;
         RECT  0.0 863.88 142.24 864.44 ;
         LAYER MET3 ;
         RECT  892.4 871.24 899.4 871.8 ;
         LAYER MET3 ;
         RECT  0.0 676.2 899.4 676.76 ;
         LAYER MET3 ;
         RECT  0.0 941.16 899.4 941.72 ;
         LAYER MET4 ;
         RECT  714.84 0.0 715.4 976.68 ;
         LAYER MET3 ;
         RECT  0.0 396.52 177.2 397.08 ;
         LAYER MET3 ;
         RECT  0.0 442.52 899.4 443.08 ;
         LAYER MET4 ;
         RECT  635.72 0.0 636.28 976.68 ;
         LAYER MET4 ;
         RECT  2.76 0.0 3.32 976.68 ;
         LAYER MET4 ;
         RECT  67.16 0.0 67.72 976.68 ;
         LAYER MET4 ;
         RECT  322.92 0.0 323.48 976.68 ;
         LAYER MET4 ;
         RECT  138.92 0.0 139.48 976.68 ;
         LAYER MET3 ;
         RECT  0.0 540.04 142.24 540.6 ;
         LAYER MET3 ;
         RECT  0.0 69.0 160.64 69.56 ;
         LAYER MET3 ;
         RECT  716.68 333.96 899.4 334.52 ;
         LAYER MET3 ;
         RECT  733.24 862.04 899.4 862.6 ;
         LAYER MET3 ;
         RECT  0.0 834.44 899.4 835.0 ;
         LAYER MET4 ;
         RECT  34.04 0.0 34.6 976.68 ;
         LAYER MET3 ;
         RECT  821.56 45.08 899.4 45.64 ;
         LAYER MET3 ;
         RECT  0.0 111.32 117.4 111.88 ;
         LAYER MET3 ;
         RECT  0.0 405.72 899.4 406.28 ;
         LAYER MET4 ;
         RECT  742.44 0.0 743.0 976.68 ;
         LAYER MET3 ;
         RECT  0.0 65.32 899.4 65.88 ;
         LAYER MET4 ;
         RECT  851.0 0.0 851.56 976.68 ;
         LAYER MET3 ;
         RECT  0.0 236.44 899.4 237.0 ;
         LAYER MET3 ;
         RECT  0.0 24.84 87.96 25.4 ;
         LAYER MET3 ;
         RECT  0.0 536.36 899.4 536.92 ;
         LAYER MET3 ;
         RECT  0.0 210.68 117.4 211.24 ;
         LAYER MET4 ;
         RECT  317.4 0.0 317.96 976.68 ;
         LAYER MET3 ;
         RECT  0.0 665.16 142.24 665.72 ;
         LAYER MET3 ;
         RECT  0.0 378.12 899.4 378.68 ;
         LAYER MET3 ;
         RECT  0.0 869.4 177.2 869.96 ;
         LAYER MET4 ;
         RECT  50.6 0.0 51.16 976.68 ;
         LAYER MET3 ;
         RECT  808.68 972.44 899.4 973.0 ;
         LAYER MET3 ;
         RECT  394.68 4.6 899.4 5.16 ;
         LAYER MET4 ;
         RECT  236.44 0.0 237.0 976.68 ;
         LAYER MET3 ;
         RECT  0.0 332.12 899.4 332.68 ;
         LAYER MET4 ;
         RECT  425.96 0.0 426.52 976.68 ;
         LAYER MET4 ;
         RECT  45.08 0.0 45.64 976.68 ;
         LAYER MET3 ;
         RECT  797.64 166.52 899.4 167.08 ;
         LAYER MET3 ;
         RECT  0.0 484.84 899.4 485.4 ;
         LAYER MET3 ;
         RECT  0.0 534.52 899.4 535.08 ;
         LAYER MET3 ;
         RECT  0.0 827.08 899.4 827.64 ;
         LAYER MET4 ;
         RECT  567.64 0.0 568.2 976.68 ;
         LAYER MET4 ;
         RECT  137.08 0.0 137.64 976.68 ;
         LAYER MET4 ;
         RECT  181.24 0.0 181.8 976.68 ;
         LAYER MET3 ;
         RECT  0.0 151.8 899.4 152.36 ;
         LAYER MET4 ;
         RECT  65.32 0.0 65.88 976.68 ;
         LAYER MET3 ;
         RECT  716.68 782.92 899.4 783.48 ;
         LAYER MET4 ;
         RECT  354.2 14.72 354.76 976.68 ;
         LAYER MET3 ;
         RECT  0.0 762.68 160.64 763.24 ;
         LAYER MET4 ;
         RECT  442.52 0.0 443.08 976.68 ;
         LAYER MET4 ;
         RECT  262.2 0.0 262.76 976.68 ;
         LAYER MET4 ;
         RECT  781.08 0.0 781.64 976.68 ;
         LAYER MET4 ;
         RECT  586.04 0.0 586.6 13.44 ;
         LAYER MET3 ;
         RECT  0.0 276.92 899.4 277.48 ;
         LAYER MET4 ;
         RECT  295.32 0.0 295.88 976.68 ;
         LAYER MET3 ;
         RECT  0.0 961.4 176.28 961.96 ;
         LAYER MET3 ;
         RECT  0.0 567.64 899.4 568.2 ;
         LAYER MET3 ;
         RECT  755.32 514.28 899.4 514.84 ;
         LAYER MET3 ;
         RECT  0.0 569.48 899.4 570.04 ;
         LAYER MET3 ;
         RECT  0.0 893.32 158.8 893.88 ;
         LAYER MET4 ;
         RECT  661.48 0.0 662.04 976.68 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER MET4 ;
         RECT  362.48 0.0 363.04 976.68 ;
         LAYER MET4 ;
         RECT  522.56 0.0 523.12 976.68 ;
         LAYER MET3 ;
         RECT  716.68 143.52 899.4 144.08 ;
         LAYER MET3 ;
         RECT  0.0 855.6 899.4 856.16 ;
         LAYER MET3 ;
         RECT  0.0 555.68 899.4 556.24 ;
         LAYER MET4 ;
         RECT  27.6 0.0 28.16 976.68 ;
         LAYER MET4 ;
         RECT  667.92 0.0 668.48 976.68 ;
         LAYER MET3 ;
         RECT  0.0 274.16 899.4 274.72 ;
         LAYER MET3 ;
         RECT  0.0 559.36 162.48 559.92 ;
         LAYER MET4 ;
         RECT  333.04 0.0 333.6 976.68 ;
         LAYER MET3 ;
         RECT  716.68 290.72 899.4 291.28 ;
         LAYER MET3 ;
         RECT  733.24 421.36 899.4 421.92 ;
         LAYER MET3 ;
         RECT  0.0 820.64 162.48 821.2 ;
         LAYER MET3 ;
         RECT  733.24 870.32 899.4 870.88 ;
         LAYER MET4 ;
         RECT  483.92 20.24 484.48 976.68 ;
         LAYER MET4 ;
         RECT  506.0 0.0 506.56 976.68 ;
         LAYER MET3 ;
         RECT  0.0 868.48 881.0 869.04 ;
         LAYER MET3 ;
         RECT  0.0 483.92 160.64 484.48 ;
         LAYER MET3 ;
         RECT  0.0 897.92 882.84 898.48 ;
         LAYER MET4 ;
         RECT  833.52 0.0 834.08 976.68 ;
         LAYER MET4 ;
         RECT  345.92 0.0 346.48 976.68 ;
         LAYER MET3 ;
         RECT  0.0 678.96 899.4 679.52 ;
         LAYER MET3 ;
         RECT  0.0 724.96 899.4 725.52 ;
         LAYER MET3 ;
         RECT  0.0 620.08 162.48 620.64 ;
         LAYER MET4 ;
         RECT  112.24 6.44 112.8 976.68 ;
         LAYER MET4 ;
         RECT  702.88 0.0 703.44 976.68 ;
         LAYER MET3 ;
         RECT  716.68 813.28 899.4 813.84 ;
         LAYER MET4 ;
         RECT  239.2 0.0 239.76 5.16 ;
         LAYER MET4 ;
         RECT  780.16 0.0 780.72 976.68 ;
         LAYER MET4 ;
         RECT  862.96 0.0 863.52 959.2 ;
         LAYER MET3 ;
         RECT  780.16 196.88 899.4 197.44 ;
         LAYER MET3 ;
         RECT  0.0 943.92 854.32 944.48 ;
         LAYER MET4 ;
         RECT  134.32 0.0 134.88 976.68 ;
         LAYER MET4 ;
         RECT  756.24 0.0 756.8 976.68 ;
         LAYER MET4 ;
         RECT  299.92 0.0 300.48 976.68 ;
         LAYER MET3 ;
         RECT  0.0 259.44 117.4 260.0 ;
         LAYER MET4 ;
         RECT  483.92 0.0 484.48 15.28 ;
         LAYER MET3 ;
         RECT  0.0 588.8 177.2 589.36 ;
         LAYER MET3 ;
         RECT  0.0 708.4 160.64 708.96 ;
         LAYER MET3 ;
         RECT  0.0 802.24 899.4 802.8 ;
         LAYER MET3 ;
         RECT  0.0 896.08 899.4 896.64 ;
         LAYER MET4 ;
         RECT  187.68 0.0 188.24 976.68 ;
         LAYER MET4 ;
         RECT  478.4 0.0 478.96 976.68 ;
         LAYER MET4 ;
         RECT  559.36 0.0 559.92 976.68 ;
         LAYER MET3 ;
         RECT  0.0 756.24 899.4 756.8 ;
         LAYER MET4 ;
         RECT  86.48 0.0 87.04 976.68 ;
         LAYER MET3 ;
         RECT  733.24 632.96 899.4 633.52 ;
         LAYER MET4 ;
         RECT  356.96 0.0 357.52 976.68 ;
         LAYER MET3 ;
         RECT  780.16 123.28 899.4 123.84 ;
         LAYER MET4 ;
         RECT  535.44 0.0 536.0 976.68 ;
         LAYER MET4 ;
         RECT  270.48 0.0 271.04 976.68 ;
         LAYER MET4 ;
         RECT  758.08 0.0 758.64 976.68 ;
         LAYER MET4 ;
         RECT  355.12 0.0 355.68 5.16 ;
         LAYER MET3 ;
         RECT  0.0 414.0 177.2 414.56 ;
         LAYER MET4 ;
         RECT  794.88 0.0 795.44 976.68 ;
         LAYER MET4 ;
         RECT  708.4 0.0 708.96 976.68 ;
         LAYER MET4 ;
         RECT  598.0 0.0 598.56 976.68 ;
         LAYER MET4 ;
         RECT  603.52 0.0 604.08 976.68 ;
         LAYER MET3 ;
         RECT  0.0 498.64 899.4 499.2 ;
         LAYER MET3 ;
         RECT  0.0 281.52 117.4 282.08 ;
         LAYER MET3 ;
         RECT  0.0 728.64 899.4 729.2 ;
         LAYER MET3 ;
         RECT  716.68 886.88 899.4 887.44 ;
         LAYER MET3 ;
         RECT  0.0 64.4 170.76 64.96 ;
         LAYER MET4 ;
         RECT  347.76 0.0 348.32 962.88 ;
         LAYER MET4 ;
         RECT  476.56 0.0 477.12 976.68 ;
         LAYER MET3 ;
         RECT  0.0 369.84 899.4 370.4 ;
         LAYER MET4 ;
         RECT  564.88 0.0 565.44 976.68 ;
         LAYER MET3 ;
         RECT  398.36 9.2 899.4 9.76 ;
         LAYER MET3 ;
         RECT  733.24 682.64 899.4 683.2 ;
         LAYER MET3 ;
         RECT  0.0 719.44 162.48 720.0 ;
         LAYER MET3 ;
         RECT  0.0 804.08 899.4 804.64 ;
         LAYER MET4 ;
         RECT  842.72 0.0 843.28 976.68 ;
         LAYER MET3 ;
         RECT  689.08 22.08 899.4 22.64 ;
         LAYER MET3 ;
         RECT  0.0 358.8 160.64 359.36 ;
         LAYER MET3 ;
         RECT  0.0 513.36 899.4 513.92 ;
         LAYER MET3 ;
         RECT  866.64 951.28 899.4 951.84 ;
         LAYER MET4 ;
         RECT  715.76 0.0 716.32 976.68 ;
         LAYER MET3 ;
         RECT  0.0 333.04 80.6 333.6 ;
         LAYER MET3 ;
         RECT  0.0 80.96 899.4 81.52 ;
         LAYER MET3 ;
         RECT  0.0 323.84 899.4 324.4 ;
         LAYER MET3 ;
         RECT  0.0 351.44 899.4 352.0 ;
         LAYER MET4 ;
         RECT  213.44 0.0 214.0 11.6 ;
         LAYER MET4 ;
         RECT  855.6 0.0 856.16 976.68 ;
         LAYER MET3 ;
         RECT  731.4 620.08 899.4 620.64 ;
         LAYER MET3 ;
         RECT  95.68 312.8 899.4 313.36 ;
         LAYER MET3 ;
         RECT  0.0 325.68 899.4 326.24 ;
         LAYER MET4 ;
         RECT  701.04 0.0 701.6 976.68 ;
         LAYER MET3 ;
         RECT  0.0 60.72 899.4 61.28 ;
         LAYER MET3 ;
         RECT  0.0 651.36 142.24 651.92 ;
         LAYER MET3 ;
         RECT  132.48 31.28 899.4 31.84 ;
         LAYER MET3 ;
         RECT  0.0 877.68 899.4 878.24 ;
         LAYER MET4 ;
         RECT  741.52 0.0 742.08 976.68 ;
         LAYER MET3 ;
         RECT  0.0 101.2 899.4 101.76 ;
         LAYER MET3 ;
         RECT  0.0 401.12 899.4 401.68 ;
         LAYER MET3 ;
         RECT  0.0 859.28 881.0 859.84 ;
         LAYER MET3 ;
         RECT  821.56 71.76 899.4 72.32 ;
         LAYER MET3 ;
         RECT  869.4 943.92 899.4 944.48 ;
         LAYER MET4 ;
         RECT  62.56 0.0 63.12 976.68 ;
         LAYER MET4 ;
         RECT  115.92 0.0 116.48 976.68 ;
         LAYER MET3 ;
         RECT  0.0 921.84 808.32 922.4 ;
         LAYER MET4 ;
         RECT  864.8 0.0 865.36 976.68 ;
         LAYER MET3 ;
         RECT  731.4 669.76 899.4 670.32 ;
         LAYER MET3 ;
         RECT  780.16 95.68 899.4 96.24 ;
         LAYER MET3 ;
         RECT  716.68 839.04 899.4 839.6 ;
         LAYER MET3 ;
         RECT  733.24 434.24 899.4 434.8 ;
         LAYER MET4 ;
         RECT  161.92 6.44 162.48 976.68 ;
         LAYER MET4 ;
         RECT  292.56 6.44 293.12 976.68 ;
         LAYER MET4 ;
         RECT  655.04 0.0 655.6 976.68 ;
         LAYER MET4 ;
         RECT  726.8 0.0 727.36 976.68 ;
         LAYER MET4 ;
         RECT  761.76 0.0 762.32 976.68 ;
         LAYER MET3 ;
         RECT  780.16 191.36 899.4 191.92 ;
         LAYER MET4 ;
         RECT  664.24 0.0 664.8 976.68 ;
         LAYER MET3 ;
         RECT  0.0 20.24 32.76 20.8 ;
         LAYER MET3 ;
         RECT  733.24 384.56 899.4 385.12 ;
         LAYER MET3 ;
         RECT  755.32 428.72 899.4 429.28 ;
         LAYER MET3 ;
         RECT  0.0 745.2 160.64 745.76 ;
         LAYER MET4 ;
         RECT  642.16 0.0 642.72 976.68 ;
         LAYER MET3 ;
         RECT  0.0 182.16 117.4 182.72 ;
         LAYER MET4 ;
         RECT  198.72 0.0 199.28 976.68 ;
         LAYER MET3 ;
         RECT  0.0 599.84 899.4 600.4 ;
         LAYER MET3 ;
         RECT  0.0 710.24 899.4 710.8 ;
         LAYER MET3 ;
         RECT  755.32 677.12 899.4 677.68 ;
         LAYER MET3 ;
         RECT  0.0 491.28 177.2 491.84 ;
         LAYER MET4 ;
         RECT  782.0 0.0 782.56 976.68 ;
         LAYER MET4 ;
         RECT  585.12 0.0 585.68 13.44 ;
         LAYER MET3 ;
         RECT  0.0 548.32 899.4 548.88 ;
         LAYER MET3 ;
         RECT  0.0 184.0 117.4 184.56 ;
         LAYER MET3 ;
         RECT  0.0 886.88 177.2 887.44 ;
         LAYER MET3 ;
         RECT  0.0 772.8 899.4 773.36 ;
         LAYER MET4 ;
         RECT  248.4 0.0 248.96 976.68 ;
         LAYER MET4 ;
         RECT  465.52 0.0 466.08 976.68 ;
         LAYER MET3 ;
         RECT  0.0 222.64 160.64 223.2 ;
         LAYER MET3 ;
         RECT  0.0 934.72 739.32 935.28 ;
         LAYER MET3 ;
         RECT  0.0 356.96 899.4 357.52 ;
         LAYER MET3 ;
         RECT  733.24 397.44 899.4 398.0 ;
         LAYER MET3 ;
         RECT  0.0 386.4 899.4 386.96 ;
         LAYER MET3 ;
         RECT  0.0 881.36 160.64 881.92 ;
         LAYER MET4 ;
         RECT  379.04 0.0 379.6 976.68 ;
         LAYER MET3 ;
         RECT  0.0 12.88 22.64 13.44 ;
         LAYER MET3 ;
         RECT  689.08 18.4 899.4 18.96 ;
         LAYER MET3 ;
         RECT  0.0 677.12 142.24 677.68 ;
         LAYER MET4 ;
         RECT  574.08 0.0 574.64 976.68 ;
         LAYER MET3 ;
         RECT  0.0 73.6 160.64 74.16 ;
         LAYER MET3 ;
         RECT  0.0 139.84 899.4 140.4 ;
         LAYER MET3 ;
         RECT  19.32 53.36 899.4 53.92 ;
         LAYER MET4 ;
         RECT  524.4 0.0 524.96 976.68 ;
         LAYER MET4 ;
         RECT  594.32 0.0 594.88 976.68 ;
         LAYER MET4 ;
         RECT  699.2 0.0 699.76 976.68 ;
         LAYER MET3 ;
         RECT  0.0 447.12 160.64 447.68 ;
         LAYER MET3 ;
         RECT  0.0 953.12 899.4 953.68 ;
         LAYER MET4 ;
         RECT  710.24 0.0 710.8 976.68 ;
         LAYER MET3 ;
         RECT  716.68 888.72 899.4 889.28 ;
         LAYER MET4 ;
         RECT  368.0 0.0 368.56 976.68 ;
         LAYER MET3 ;
         RECT  0.0 209.76 117.4 210.32 ;
         LAYER MET4 ;
         RECT  136.16 0.0 136.72 976.68 ;
         LAYER MET3 ;
         RECT  0.0 93.84 117.4 94.4 ;
         LAYER MET3 ;
         RECT  0.0 172.96 117.4 173.52 ;
         LAYER MET3 ;
         RECT  0.0 390.08 177.2 390.64 ;
         LAYER MET3 ;
         RECT  0.0 798.56 899.4 799.12 ;
         LAYER MET3 ;
         RECT  0.0 844.56 160.64 845.12 ;
         LAYER MET3 ;
         RECT  0.0 195.04 117.4 195.6 ;
         LAYER MET3 ;
         RECT  0.0 885.04 881.0 885.6 ;
         LAYER MET3 ;
         RECT  0.0 480.24 899.4 480.8 ;
         LAYER MET3 ;
         RECT  0.0 750.72 142.24 751.28 ;
         LAYER MET3 ;
         RECT  0.0 971.52 752.2 972.08 ;
         LAYER MET4 ;
         RECT  586.96 0.0 587.52 976.68 ;
         LAYER MET3 ;
         RECT  0.0 196.88 117.4 197.44 ;
         LAYER MET3 ;
         RECT  0.0 826.16 142.24 826.72 ;
         LAYER MET3 ;
         RECT  0.0 314.64 177.2 315.2 ;
         LAYER MET4 ;
         RECT  754.4 0.0 754.96 970.24 ;
         LAYER MET4 ;
         RECT  402.96 0.0 403.52 976.68 ;
         LAYER MET3 ;
         RECT  0.0 257.6 117.4 258.16 ;
         LAYER MET4 ;
         RECT  485.76 0.0 486.32 976.68 ;
         LAYER MET3 ;
         RECT  0.0 916.32 179.04 916.88 ;
         LAYER MET4 ;
         RECT  163.76 0.0 164.32 976.68 ;
         LAYER MET3 ;
         RECT  0.0 958.64 860.76 959.2 ;
         LAYER MET3 ;
         RECT  0.0 494.96 899.4 495.52 ;
         LAYER MET3 ;
         RECT  733.24 198.72 899.4 199.28 ;
         LAYER MET3 ;
         RECT  96.6 320.16 899.4 320.72 ;
         LAYER MET3 ;
         RECT  0.0 5.52 110.04 6.08 ;
         LAYER MET4 ;
         RECT  421.36 0.0 421.92 976.68 ;
         LAYER MET3 ;
         RECT  0.0 695.52 160.64 696.08 ;
         LAYER MET3 ;
         RECT  0.0 522.56 899.4 523.12 ;
         LAYER MET3 ;
         RECT  0.0 662.4 899.4 662.96 ;
         LAYER MET4 ;
         RECT  84.64 0.0 85.2 976.68 ;
         LAYER MET4 ;
         RECT  778.32 0.0 778.88 976.68 ;
         LAYER MET3 ;
         RECT  780.16 285.2 899.4 285.76 ;
         LAYER MET3 ;
         RECT  716.68 391.92 899.4 392.48 ;
         LAYER MET3 ;
         RECT  0.0 268.64 117.4 269.2 ;
         LAYER MET4 ;
         RECT  158.24 0.0 158.8 976.68 ;
         LAYER MET4 ;
         RECT  51.52 0.0 52.08 976.68 ;
         LAYER MET3 ;
         RECT  780.16 132.48 899.4 133.04 ;
         LAYER MET3 ;
         RECT  0.0 920.0 899.4 920.56 ;
         LAYER MET3 ;
         RECT  780.16 281.52 899.4 282.08 ;
         LAYER MET3 ;
         RECT  0.0 853.76 899.4 854.32 ;
         LAYER MET3 ;
         RECT  0.0 969.68 899.4 970.24 ;
         LAYER MET3 ;
         RECT  0.0 362.48 899.4 363.04 ;
         LAYER MET3 ;
         RECT  0.0 629.28 899.4 629.84 ;
         LAYER MET3 ;
         RECT  821.56 55.2 899.4 55.76 ;
         LAYER MET3 ;
         RECT  868.48 964.16 899.4 964.72 ;
         LAYER MET4 ;
         RECT  11.04 0.0 11.6 976.68 ;
         LAYER MET4 ;
         RECT  800.4 0.0 800.96 976.68 ;
         LAYER MET3 ;
         RECT  0.0 789.36 177.2 789.92 ;
         LAYER MET3 ;
         RECT  0.0 666.08 899.4 666.64 ;
         LAYER MET3 ;
         RECT  0.0 903.44 899.4 904.0 ;
         LAYER MET3 ;
         RECT  0.0 581.44 899.4 582.0 ;
         LAYER MET4 ;
         RECT  375.36 0.0 375.92 976.68 ;
         LAYER MET3 ;
         RECT  0.0 288.88 899.4 289.44 ;
         LAYER MET3 ;
         RECT  0.0 474.72 899.4 475.28 ;
         LAYER MET3 ;
         RECT  0.0 165.6 177.2 166.16 ;
         LAYER MET3 ;
         RECT  821.56 79.12 899.4 79.68 ;
         LAYER MET3 ;
         RECT  780.16 242.88 899.4 243.44 ;
         LAYER MET4 ;
         RECT  494.96 0.0 495.52 976.68 ;
         LAYER MET3 ;
         RECT  0.0 669.76 162.48 670.32 ;
         LAYER MET4 ;
         RECT  504.16 0.0 504.72 976.68 ;
         LAYER MET3 ;
         RECT  0.0 276.0 899.4 276.56 ;
         LAYER MET3 ;
         RECT  83.72 299.92 899.4 300.48 ;
         LAYER MET3 ;
         RECT  0.0 342.24 177.2 342.8 ;
         LAYER MET4 ;
         RECT  180.32 20.24 180.88 976.68 ;
         LAYER MET3 ;
         RECT  0.0 458.16 162.48 458.72 ;
         LAYER MET4 ;
         RECT  460.0 0.0 460.56 976.68 ;
         LAYER MET3 ;
         RECT  733.24 831.68 899.4 832.24 ;
         LAYER MET3 ;
         RECT  733.24 248.4 899.4 248.96 ;
         LAYER MET4 ;
         RECT  145.36 0.0 145.92 976.68 ;
         LAYER MET3 ;
         RECT  0.0 242.88 117.4 243.44 ;
         LAYER MET4 ;
         RECT  322.0 0.0 322.56 5.16 ;
         LAYER MET4 ;
         RECT  338.56 18.4 339.12 976.68 ;
         LAYER MET4 ;
         RECT  706.56 0.0 707.12 976.68 ;
         LAYER MET3 ;
         RECT  0.0 504.16 899.4 504.72 ;
         LAYER MET3 ;
         RECT  0.0 18.4 30.0 18.96 ;
         LAYER MET3 ;
         RECT  0.0 862.96 177.2 863.52 ;
         LAYER MET3 ;
         RECT  0.0 292.56 177.2 293.12 ;
         LAYER MET3 ;
         RECT  0.0 279.68 100.84 280.24 ;
         LAYER MET4 ;
         RECT  123.28 0.0 123.84 976.68 ;
         LAYER MET4 ;
         RECT  404.8 0.0 405.36 5.16 ;
         LAYER MET3 ;
         RECT  780.16 180.32 899.4 180.88 ;
         LAYER MET4 ;
         RECT  743.36 0.0 743.92 976.68 ;
         LAYER MET3 ;
         RECT  0.0 187.68 899.4 188.24 ;
         LAYER MET4 ;
         RECT  404.8 20.24 405.36 976.68 ;
         LAYER MET4 ;
         RECT  599.84 0.0 600.4 976.68 ;
         LAYER MET4 ;
         RECT  879.52 0.0 880.08 976.68 ;
         LAYER MET3 ;
         RECT  755.32 228.16 899.4 228.72 ;
         LAYER MET3 ;
         RECT  780.16 270.48 899.4 271.04 ;
         LAYER MET3 ;
         RECT  0.0 294.4 73.24 294.96 ;
         LAYER MET4 ;
         RECT  314.64 0.0 315.2 11.6 ;
         LAYER MET3 ;
         RECT  755.32 353.28 899.4 353.84 ;
         LAYER MET4 ;
         RECT  719.44 0.0 720.0 976.68 ;
         LAYER MET3 ;
         RECT  0.0 382.72 899.4 383.28 ;
         LAYER MET4 ;
         RECT  309.12 0.0 309.68 976.68 ;
         LAYER MET4 ;
         RECT  820.64 71.76 821.2 976.68 ;
         LAYER MET4 ;
         RECT  866.64 0.0 867.2 976.68 ;
         LAYER MET3 ;
         RECT  0.0 634.8 899.4 635.36 ;
         LAYER MET3 ;
         RECT  0.0 759.92 899.4 760.48 ;
         LAYER MET4 ;
         RECT  563.04 0.0 563.6 976.68 ;
         LAYER MET3 ;
         RECT  0.0 540.96 177.2 541.52 ;
         LAYER MET4 ;
         RECT  180.32 0.0 180.88 9.76 ;
         LAYER MET3 ;
         RECT  0.0 496.8 160.64 497.36 ;
         LAYER MET4 ;
         RECT  288.88 0.0 289.44 5.16 ;
         LAYER MET3 ;
         RECT  780.16 266.8 899.4 267.36 ;
         LAYER MET3 ;
         RECT  91.08 33.12 899.4 33.68 ;
         LAYER MET4 ;
         RECT  143.52 6.44 144.08 976.68 ;
         LAYER MET3 ;
         RECT  0.0 143.52 177.2 144.08 ;
         LAYER MET4 ;
         RECT  323.84 0.0 324.4 976.68 ;
         LAYER MET4 ;
         RECT  426.88 0.0 427.44 976.68 ;
         LAYER MET3 ;
         RECT  733.24 583.28 899.4 583.84 ;
         LAYER MET4 ;
         RECT  154.56 0.0 155.12 976.68 ;
         LAYER MET3 ;
         RECT  0.0 329.36 77.84 329.92 ;
         LAYER MET3 ;
         RECT  733.24 358.8 899.4 359.36 ;
         LAYER MET4 ;
         RECT  653.2 0.0 653.76 9.76 ;
         LAYER MET4 ;
         RECT  12.88 0.0 13.44 976.68 ;
         LAYER MET4 ;
         RECT  75.44 0.0 76.0 976.68 ;
         LAYER MET3 ;
         RECT  0.0 726.8 142.24 727.36 ;
         LAYER MET3 ;
         RECT  0.0 327.52 899.4 328.08 ;
         LAYER MET4 ;
         RECT  58.88 0.0 59.44 976.68 ;
         LAYER MET3 ;
         RECT  17.48 42.32 899.4 42.88 ;
         LAYER MET3 ;
         RECT  0.0 128.8 100.84 129.36 ;
         LAYER MET3 ;
         RECT  0.0 316.48 80.6 317.04 ;
         LAYER MET3 ;
         RECT  0.0 636.64 899.4 637.2 ;
         LAYER MET4 ;
         RECT  316.48 0.0 317.04 976.68 ;
         LAYER MET4 ;
         RECT  342.24 6.44 342.8 976.68 ;
         LAYER MET4 ;
         RECT  572.24 0.0 572.8 976.68 ;
         LAYER MET3 ;
         RECT  0.0 395.6 899.4 396.16 ;
         LAYER MET3 ;
         RECT  17.48 75.44 899.4 76.0 ;
         LAYER MET4 ;
         RECT  303.6 0.0 304.16 976.68 ;
         LAYER MET4 ;
         RECT  815.12 0.0 815.68 976.68 ;
         LAYER MET4 ;
         RECT  724.96 0.0 725.52 976.68 ;
         LAYER MET4 ;
         RECT  739.68 0.0 740.24 976.68 ;
         LAYER MET3 ;
         RECT  0.0 49.68 87.96 50.24 ;
         LAYER MET3 ;
         RECT  0.0 842.72 899.4 843.28 ;
         LAYER MET4 ;
         RECT  263.12 0.0 263.68 976.68 ;
         LAYER MET3 ;
         RECT  0.0 951.28 766.0 951.84 ;
         LAYER MET3 ;
         RECT  0.0 68.08 815.68 68.64 ;
         LAYER MET3 ;
         RECT  826.16 90.16 899.4 90.72 ;
         LAYER MET4 ;
         RECT  874.0 0.0 874.56 976.68 ;
         LAYER MET3 ;
         RECT  0.0 228.16 142.24 228.72 ;
         LAYER MET3 ;
         RECT  0.0 11.04 5.16 11.6 ;
         LAYER MET3 ;
         RECT  755.32 651.36 899.4 651.92 ;
         LAYER MET3 ;
         RECT  0.0 691.84 899.4 692.4 ;
         LAYER MET3 ;
         RECT  797.64 204.24 899.4 204.8 ;
         LAYER MET3 ;
         RECT  0.0 787.52 177.2 788.08 ;
         LAYER MET3 ;
         RECT  0.0 758.08 160.64 758.64 ;
         LAYER MET3 ;
         RECT  0.0 918.16 752.2 918.72 ;
         LAYER MET4 ;
         RECT  837.2 0.0 837.76 976.68 ;
         LAYER MET4 ;
         RECT  125.12 0.0 125.68 976.68 ;
         LAYER MET3 ;
         RECT  0.0 701.04 142.24 701.6 ;
         LAYER MET4 ;
         RECT  434.24 0.0 434.8 976.68 ;
         LAYER MET3 ;
         RECT  0.0 167.44 117.4 168.0 ;
         LAYER MET3 ;
         RECT  0.0 174.8 899.4 175.36 ;
         LAYER MET3 ;
         RECT  0.0 872.16 899.4 872.72 ;
         LAYER MET4 ;
         RECT  653.2 20.24 653.76 976.68 ;
         LAYER MET4 ;
         RECT  861.12 0.0 861.68 959.2 ;
         LAYER MET3 ;
         RECT  0.0 645.84 160.64 646.4 ;
         LAYER MET3 ;
         RECT  0.0 851.92 899.4 852.48 ;
         LAYER MET3 ;
         RECT  780.16 169.28 899.4 169.84 ;
         LAYER MET4 ;
         RECT  349.6 20.24 350.16 976.68 ;
         LAYER MET4 ;
         RECT  310.96 6.44 311.52 976.68 ;
         LAYER MET4 ;
         RECT  811.44 0.0 812.0 976.68 ;
         LAYER MET3 ;
         RECT  780.16 184.0 899.4 184.56 ;
         LAYER MET4 ;
         RECT  491.28 0.0 491.84 976.68 ;
         LAYER MET3 ;
         RECT  0.0 189.52 899.4 190.08 ;
         LAYER MET3 ;
         RECT  716.68 540.96 899.4 541.52 ;
         LAYER MET3 ;
         RECT  0.0 828.0 899.4 828.56 ;
         LAYER MET4 ;
         RECT  447.12 0.0 447.68 962.88 ;
         LAYER MET3 ;
         RECT  0.0 104.88 100.84 105.44 ;
         LAYER MET3 ;
         RECT  0.0 334.88 160.64 335.44 ;
         LAYER MET4 ;
         RECT  425.04 0.0 425.6 976.68 ;
         LAYER MET3 ;
         RECT  0.0 412.16 899.4 412.72 ;
         LAYER MET4 ;
         RECT  540.96 0.0 541.52 976.68 ;
         LAYER MET4 ;
         RECT  769.12 0.0 769.68 970.24 ;
         LAYER MET3 ;
         RECT  0.0 938.4 808.32 938.96 ;
         LAYER MET3 ;
         RECT  755.32 826.16 899.4 826.72 ;
         LAYER MET4 ;
         RECT  783.84 0.0 784.4 976.68 ;
         LAYER MET3 ;
         RECT  755.32 601.68 899.4 602.24 ;
         LAYER MET3 ;
         RECT  0.0 537.28 899.4 537.84 ;
         LAYER MET4 ;
         RECT  182.16 0.0 182.72 976.68 ;
         LAYER MET3 ;
         RECT  0.0 126.96 899.4 127.52 ;
         LAYER MET3 ;
         RECT  0.0 482.08 899.4 482.64 ;
         LAYER MET4 ;
         RECT  314.64 20.24 315.2 976.68 ;
         LAYER MET4 ;
         RECT  736.0 0.0 736.56 976.68 ;
         LAYER MET3 ;
         RECT  780.16 108.56 899.4 109.12 ;
         LAYER MET4 ;
         RECT  437.92 0.0 438.48 976.68 ;
         LAYER MET4 ;
         RECT  544.64 0.0 545.2 976.68 ;
         LAYER MET3 ;
         RECT  733.24 471.04 899.4 471.6 ;
         LAYER MET3 ;
         RECT  0.0 612.72 899.4 613.28 ;
         LAYER MET4 ;
         RECT  121.44 0.0 122.0 976.68 ;
         LAYER MET3 ;
         RECT  0.0 309.12 160.64 309.68 ;
         LAYER MET3 ;
         RECT  716.68 115.92 899.4 116.48 ;
         LAYER MET4 ;
         RECT  487.6 0.0 488.16 976.68 ;
         LAYER MET4 ;
         RECT  305.44 0.0 306.0 5.16 ;
         LAYER MET4 ;
         RECT  207.92 0.0 208.48 976.68 ;
         LAYER MET3 ;
         RECT  0.0 84.64 815.68 85.2 ;
         LAYER MET4 ;
         RECT  688.16 0.0 688.72 17.12 ;
         LAYER MET3 ;
         RECT  0.0 644.0 899.4 644.56 ;
         LAYER MET4 ;
         RECT  419.52 0.0 420.08 976.68 ;
         LAYER MET4 ;
         RECT  47.84 0.0 48.4 976.68 ;
         LAYER MET4 ;
         RECT  224.48 0.0 225.04 976.68 ;
         LAYER MET4 ;
         RECT  579.6 0.0 580.16 976.68 ;
         LAYER MET4 ;
         RECT  93.84 0.0 94.4 976.68 ;
         LAYER MET4 ;
         RECT  680.8 0.0 681.36 976.68 ;
         LAYER MET4 ;
         RECT  840.88 0.0 841.44 976.68 ;
         LAYER MET4 ;
         RECT  97.52 0.0 98.08 976.68 ;
         LAYER MET4 ;
         RECT  95.68 0.0 96.24 976.68 ;
         LAYER MET3 ;
         RECT  780.16 106.72 899.4 107.28 ;
         LAYER MET4 ;
         RECT  388.24 12.88 388.8 976.68 ;
         LAYER MET3 ;
         RECT  80.04 310.96 899.4 311.52 ;
         LAYER MET3 ;
         RECT  0.0 945.76 899.4 946.32 ;
         LAYER MET3 ;
         RECT  0.0 456.32 899.4 456.88 ;
         LAYER MET3 ;
         RECT  0.0 193.2 117.4 193.76 ;
         LAYER MET4 ;
         RECT  366.16 0.0 366.72 976.68 ;
         LAYER MET3 ;
         RECT  733.24 520.72 899.4 521.28 ;
         LAYER MET3 ;
         RECT  0.0 815.12 177.2 815.68 ;
         LAYER MET3 ;
         RECT  0.0 706.56 899.4 707.12 ;
         LAYER MET3 ;
         RECT  0.0 161.92 899.4 162.48 ;
         LAYER MET4 ;
         RECT  493.12 0.0 493.68 976.68 ;
         LAYER MET3 ;
         RECT  0.0 850.08 142.24 850.64 ;
         LAYER MET4 ;
         RECT  896.08 0.0 896.64 976.68 ;
         LAYER MET3 ;
         RECT  0.0 627.44 142.24 628.0 ;
         LAYER MET4 ;
         RECT  399.28 0.0 399.84 976.68 ;
         LAYER MET4 ;
         RECT  22.08 0.0 22.64 976.68 ;
         LAYER MET3 ;
         RECT  0.0 542.8 899.4 543.36 ;
         LAYER MET4 ;
         RECT  509.68 0.0 510.24 976.68 ;
         LAYER MET4 ;
         RECT  553.84 0.0 554.4 976.68 ;
         LAYER MET4 ;
         RECT  730.48 0.0 731.04 976.68 ;
         LAYER MET3 ;
         RECT  0.0 601.68 142.24 602.24 ;
         LAYER MET3 ;
         RECT  38.64 51.52 899.4 52.08 ;
         LAYER MET3 ;
         RECT  0.0 239.2 899.4 239.76 ;
         LAYER MET3 ;
         RECT  797.64 128.8 899.4 129.36 ;
         LAYER MET3 ;
         RECT  716.68 340.4 899.4 340.96 ;
         LAYER MET4 ;
         RECT  215.28 0.0 215.84 976.68 ;
         LAYER MET3 ;
         RECT  0.0 57.04 899.4 57.6 ;
         LAYER MET3 ;
         RECT  780.16 97.52 899.4 98.08 ;
         LAYER MET3 ;
         RECT  0.0 9.2 31.84 9.76 ;
         LAYER MET3 ;
         RECT  0.0 487.6 899.4 488.16 ;
         LAYER MET4 ;
         RECT  90.16 0.0 90.72 976.68 ;
         LAYER MET4 ;
         RECT  206.08 14.72 206.64 976.68 ;
         LAYER MET3 ;
         RECT  0.0 347.76 160.64 348.32 ;
         LAYER MET3 ;
         RECT  0.0 697.36 899.4 697.92 ;
         LAYER MET3 ;
         RECT  0.0 813.28 177.2 813.84 ;
         LAYER MET4 ;
         RECT  241.04 0.0 241.6 976.68 ;
         LAYER MET4 ;
         RECT  666.08 0.0 666.64 976.68 ;
         LAYER MET3 ;
         RECT  731.4 458.16 899.4 458.72 ;
         LAYER MET3 ;
         RECT  0.0 277.84 899.4 278.4 ;
         LAYER MET3 ;
         RECT  731.4 609.04 899.4 609.6 ;
         LAYER MET3 ;
         RECT  731.4 719.44 899.4 720.0 ;
         LAYER MET3 ;
         RECT  0.0 371.68 160.64 372.24 ;
         LAYER MET3 ;
         RECT  0.0 879.52 899.4 880.08 ;
         LAYER MET3 ;
         RECT  405.72 3.68 899.4 4.24 ;
         LAYER MET3 ;
         RECT  733.24 309.12 899.4 309.68 ;
         LAYER MET3 ;
         RECT  0.0 430.56 899.4 431.12 ;
         LAYER MET4 ;
         RECT  371.68 0.0 372.24 5.16 ;
         LAYER MET4 ;
         RECT  515.2 0.0 515.76 976.68 ;
         LAYER MET3 ;
         RECT  0.0 914.48 882.84 915.04 ;
         LAYER MET3 ;
         RECT  0.0 114.08 899.4 114.64 ;
         LAYER MET4 ;
         RECT  518.88 0.0 519.44 11.6 ;
         LAYER MET4 ;
         RECT  71.76 0.0 72.32 976.68 ;
         LAYER MET3 ;
         RECT  0.0 640.32 177.2 640.88 ;
         LAYER MET4 ;
         RECT  647.68 0.0 648.24 976.68 ;
         LAYER MET4 ;
         RECT  712.08 0.0 712.64 976.68 ;
         LAYER MET4 ;
         RECT  767.28 0.0 767.84 976.68 ;
         LAYER MET3 ;
         RECT  0.0 176.64 899.4 177.2 ;
         LAYER MET3 ;
         RECT  797.64 279.68 899.4 280.24 ;
         LAYER MET3 ;
         RECT  0.0 441.6 177.2 442.16 ;
         LAYER MET4 ;
         RECT  612.72 0.0 613.28 976.68 ;
         LAYER MET3 ;
         RECT  755.32 502.32 899.4 502.88 ;
         LAYER MET4 ;
         RECT  531.76 0.0 532.32 976.68 ;
         LAYER MET4 ;
         RECT  601.68 0.0 602.24 976.68 ;
         LAYER MET3 ;
         RECT  0.0 115.92 177.2 116.48 ;
         LAYER MET3 ;
         RECT  19.32 69.92 899.4 70.48 ;
         LAYER MET3 ;
         RECT  716.68 815.12 899.4 815.68 ;
         LAYER MET3 ;
         RECT  0.0 202.4 899.4 202.96 ;
         LAYER MET3 ;
         RECT  0.0 253.92 100.84 254.48 ;
         LAYER MET3 ;
         RECT  0.0 421.36 160.64 421.92 ;
         LAYER MET4 ;
         RECT  204.24 0.0 204.8 976.68 ;
         LAYER MET4 ;
         RECT  607.2 0.0 607.76 976.68 ;
         LAYER MET4 ;
         RECT  432.4 0.0 432.96 976.68 ;
         LAYER MET3 ;
         RECT  0.0 579.6 899.4 580.16 ;
         LAYER MET3 ;
         RECT  0.0 27.6 30.92 28.16 ;
         LAYER MET4 ;
         RECT  618.24 0.0 618.8 976.68 ;
         LAYER MET4 ;
         RECT  645.84 0.0 646.4 976.68 ;
         LAYER MET3 ;
         RECT  0.0 264.96 177.2 265.52 ;
         LAYER MET3 ;
         RECT  731.4 509.68 899.4 510.24 ;
         LAYER MET4 ;
         RECT  117.76 0.0 118.32 976.68 ;
         LAYER MET4 ;
         RECT  276.0 6.44 276.56 976.68 ;
         LAYER MET3 ;
         RECT  0.0 263.12 899.4 263.68 ;
         LAYER MET3 ;
         RECT  892.4 862.96 899.4 863.52 ;
         LAYER MET4 ;
         RECT  277.84 0.0 278.4 962.88 ;
         LAYER MET3 ;
         RECT  158.24 38.64 899.4 39.2 ;
         LAYER MET3 ;
         RECT  780.16 272.32 899.4 272.88 ;
         LAYER MET4 ;
         RECT  218.96 0.0 219.52 976.68 ;
         LAYER MET4 ;
         RECT  351.44 0.0 352.0 976.68 ;
         LAYER MET3 ;
         RECT  780.16 92.0 899.4 92.56 ;
         LAYER MET3 ;
         RECT  733.24 73.6 899.4 74.16 ;
         LAYER MET3 ;
         RECT  0.0 515.2 177.2 515.76 ;
         LAYER MET3 ;
         RECT  755.32 402.96 899.4 403.52 ;
         LAYER MET4 ;
         RECT  373.52 0.0 374.08 976.68 ;
         LAYER MET4 ;
         RECT  828.0 0.0 828.56 976.68 ;
         LAYER MET3 ;
         RECT  0.0 664.24 899.4 664.8 ;
         LAYER MET4 ;
         RECT  283.36 0.0 283.92 976.68 ;
         LAYER MET3 ;
         RECT  733.24 894.24 899.4 894.8 ;
         LAYER MET3 ;
         RECT  0.0 443.44 899.4 444.0 ;
         LAYER MET3 ;
         RECT  892.4 914.48 899.4 915.04 ;
         LAYER MET3 ;
         RECT  0.0 178.48 100.84 179.04 ;
         LAYER MET4 ;
         RECT  364.32 0.0 364.88 976.68 ;
         LAYER MET4 ;
         RECT  537.28 0.0 537.84 976.68 ;
         LAYER MET3 ;
         RECT  0.0 811.44 899.4 812.0 ;
         LAYER MET4 ;
         RECT  73.6 0.0 74.16 976.68 ;
         LAYER MET4 ;
         RECT  539.12 0.0 539.68 976.68 ;
         LAYER MET3 ;
         RECT  0.0 200.56 899.4 201.12 ;
         LAYER MET3 ;
         RECT  0.0 82.8 899.4 83.36 ;
         LAYER MET3 ;
         RECT  0.0 88.32 142.24 88.88 ;
         LAYER MET3 ;
         RECT  780.16 244.72 899.4 245.28 ;
         LAYER MET3 ;
         RECT  0.0 739.68 177.2 740.24 ;
         LAYER MET3 ;
         RECT  0.0 355.12 899.4 355.68 ;
         LAYER MET3 ;
         RECT  0.0 947.6 899.4 948.16 ;
         LAYER MET4 ;
         RECT  868.48 0.0 869.04 976.68 ;
         LAYER MET4 ;
         RECT  848.24 0.0 848.8 976.68 ;
         LAYER MET3 ;
         RECT  0.0 71.76 802.8 72.32 ;
         LAYER MET3 ;
         RECT  780.16 261.28 899.4 261.84 ;
         LAYER MET3 ;
         RECT  0.0 423.2 899.4 423.76 ;
         LAYER MET4 ;
         RECT  20.24 0.0 20.8 976.68 ;
         LAYER MET3 ;
         RECT  0.0 399.28 899.4 399.84 ;
         LAYER MET3 ;
         RECT  714.84 64.4 899.4 64.96 ;
         LAYER MET3 ;
         RECT  655.04 11.04 899.4 11.6 ;
         LAYER MET4 ;
         RECT  322.0 12.88 322.56 976.68 ;
         LAYER MET3 ;
         RECT  0.0 1.84 899.4 2.4 ;
         LAYER MET3 ;
         RECT  0.0 936.56 899.4 937.12 ;
         LAYER MET4 ;
         RECT  334.88 0.0 335.44 976.68 ;
         LAYER MET4 ;
         RECT  285.2 0.0 285.76 976.68 ;
         LAYER MET4 ;
         RECT  165.6 0.0 166.16 976.68 ;
         LAYER MET4 ;
         RECT  305.44 16.56 306.0 976.68 ;
         LAYER MET4 ;
         RECT  380.88 0.0 381.44 962.88 ;
         LAYER MET3 ;
         RECT  0.0 737.84 177.2 738.4 ;
         LAYER MET3 ;
         RECT  0.0 535.44 899.4 536.0 ;
         LAYER MET3 ;
         RECT  0.0 380.88 899.4 381.44 ;
         LAYER MET3 ;
         RECT  716.68 390.08 899.4 390.64 ;
         LAYER MET4 ;
         RECT  640.32 0.0 640.88 976.68 ;
         LAYER MET4 ;
         RECT  517.04 0.0 517.6 962.88 ;
         LAYER MET3 ;
         RECT  733.24 807.76 899.4 808.32 ;
         LAYER MET4 ;
         RECT  772.8 0.0 773.36 976.68 ;
         LAYER MET4 ;
         RECT  804.08 0.0 804.64 976.68 ;
         LAYER MET3 ;
         RECT  0.0 261.28 117.4 261.84 ;
         LAYER MET3 ;
         RECT  0.0 778.32 899.4 778.88 ;
         LAYER MET3 ;
         RECT  0.0 575.92 899.4 576.48 ;
         LAYER MET3 ;
         RECT  0.0 973.36 741.16 973.92 ;
         LAYER MET3 ;
         RECT  780.16 259.44 899.4 260.0 ;
         LAYER MET3 ;
         RECT  0.0 448.96 899.4 449.52 ;
         LAYER MET3 ;
         RECT  821.56 46.0 899.4 46.56 ;
         LAYER MET3 ;
         RECT  0.0 108.56 7.0 109.12 ;
         LAYER MET3 ;
         RECT  0.0 465.52 177.2 466.08 ;
         LAYER MET4 ;
         RECT  80.96 0.0 81.52 976.68 ;
         LAYER MET4 ;
         RECT  807.76 0.0 808.32 976.68 ;
         LAYER MET3 ;
         RECT  716.68 292.56 899.4 293.12 ;
         LAYER MET4 ;
         RECT  430.56 0.0 431.12 976.68 ;
         LAYER MET3 ;
         RECT  0.0 761.76 899.4 762.32 ;
         LAYER MET4 ;
         RECT  745.2 0.0 745.76 976.68 ;
         LAYER MET3 ;
         RECT  733.24 533.6 899.4 534.16 ;
         LAYER MET3 ;
         RECT  0.0 250.24 899.4 250.8 ;
         LAYER MET4 ;
         RECT  252.08 0.0 252.64 976.68 ;
         LAYER MET3 ;
         RECT  0.0 767.28 899.4 767.84 ;
         LAYER MET4 ;
         RECT  662.4 0.0 662.96 976.68 ;
         LAYER MET3 ;
         RECT  780.16 93.84 899.4 94.4 ;
         LAYER MET3 ;
         RECT  0.0 338.56 899.4 339.12 ;
         LAYER MET3 ;
         RECT  0.0 511.52 899.4 512.08 ;
         LAYER MET4 ;
         RECT  149.04 0.0 149.6 976.68 ;
         LAYER MET4 ;
         RECT  629.28 0.0 629.84 976.68 ;
         LAYER MET3 ;
         RECT  0.0 213.44 899.4 214.0 ;
         LAYER MET4 ;
         RECT  132.48 0.0 133.04 976.68 ;
         LAYER MET3 ;
         RECT  0.0 373.52 899.4 374.08 ;
         LAYER MET4 ;
         RECT  325.68 0.0 326.24 976.68 ;
         LAYER MET4 ;
         RECT  507.84 0.0 508.4 976.68 ;
         LAYER MET3 ;
         RECT  0.0 533.6 160.64 534.16 ;
         LAYER MET3 ;
         RECT  0.0 899.76 753.12 900.32 ;
         LAYER MET3 ;
         RECT  0.0 574.08 899.4 574.64 ;
         LAYER MET3 ;
         RECT  0.0 154.56 142.24 155.12 ;
         LAYER MET4 ;
         RECT  897.92 0.0 898.48 858.92 ;
         LAYER MET3 ;
         RECT  0.0 163.76 899.4 164.32 ;
         LAYER MET4 ;
         RECT  110.4 0.0 110.96 976.68 ;
         LAYER MET3 ;
         RECT  733.24 758.08 899.4 758.64 ;
         LAYER MET4 ;
         RECT  25.76 0.0 26.32 976.68 ;
         LAYER MET3 ;
         RECT  0.0 949.44 899.4 950.0 ;
         LAYER MET4 ;
         RECT  482.08 0.0 482.64 962.88 ;
         LAYER MET4 ;
         RECT  253.92 0.0 254.48 976.68 ;
         LAYER MET4 ;
         RECT  550.16 0.0 550.72 962.88 ;
         LAYER MET3 ;
         RECT  0.0 748.88 899.4 749.44 ;
         LAYER MET4 ;
         RECT  634.8 0.0 635.36 976.68 ;
         LAYER MET4 ;
         RECT  542.8 0.0 543.36 976.68 ;
         LAYER MET4 ;
         RECT  336.72 0.0 337.28 976.68 ;
         LAYER MET3 ;
         RECT  0.0 623.76 899.4 624.32 ;
         LAYER MET3 ;
         RECT  797.64 104.88 899.4 105.44 ;
         LAYER MET3 ;
         RECT  809.6 927.36 899.4 927.92 ;
         LAYER MET3 ;
         RECT  892.4 931.04 899.4 931.6 ;
         LAYER MET4 ;
         RECT  397.44 0.0 398.0 976.68 ;
         LAYER MET3 ;
         RECT  0.0 839.04 177.2 839.6 ;
         LAYER MET3 ;
         RECT  780.16 255.76 899.4 256.32 ;
         LAYER MET4 ;
         RECT  150.88 0.0 151.44 976.68 ;
         LAYER MET4 ;
         RECT  353.28 0.0 353.84 976.68 ;
         LAYER MET3 ;
         RECT  0.0 835.36 899.4 835.92 ;
         LAYER MET3 ;
         RECT  0.0 592.48 899.4 593.04 ;
         LAYER MET4 ;
         RECT  272.32 16.56 272.88 976.68 ;
         LAYER MET3 ;
         RECT  0.0 36.8 899.4 37.36 ;
         LAYER MET3 ;
         RECT  0.0 301.76 899.4 302.32 ;
         LAYER MET3 ;
         RECT  0.0 553.84 899.4 554.4 ;
         LAYER MET3 ;
         RECT  0.0 829.84 899.4 830.4 ;
         LAYER MET3 ;
         RECT  0.0 910.8 899.4 911.36 ;
         LAYER MET4 ;
         RECT  677.12 0.0 677.68 976.68 ;
         LAYER MET3 ;
         RECT  780.16 167.44 899.4 168.0 ;
         LAYER MET3 ;
         RECT  768.2 966.0 899.4 966.56 ;
         LAYER MET3 ;
         RECT  0.0 14.72 271.04 15.28 ;
         LAYER MET3 ;
         RECT  0.0 244.72 117.4 245.28 ;
         LAYER MET3 ;
         RECT  821.56 62.56 899.4 63.12 ;
         LAYER MET3 ;
         RECT  0.0 864.8 177.2 865.36 ;
         LAYER MET3 ;
         RECT  0.0 732.32 160.64 732.88 ;
         LAYER MET4 ;
         RECT  415.84 0.0 416.4 13.44 ;
         LAYER MET3 ;
         RECT  0.0 603.52 899.4 604.08 ;
         LAYER MET3 ;
         RECT  0.0 785.68 899.4 786.24 ;
         LAYER MET3 ;
         RECT  0.0 415.84 177.2 416.4 ;
         LAYER MET3 ;
         RECT  0.0 752.56 899.4 753.12 ;
         LAYER MET3 ;
         RECT  755.32 800.4 899.4 800.96 ;
         LAYER MET4 ;
         RECT  31.28 0.0 31.84 976.68 ;
         LAYER MET4 ;
         RECT  776.48 0.0 777.04 976.68 ;
         LAYER MET4 ;
         RECT  886.88 0.0 887.44 976.68 ;
         LAYER MET3 ;
         RECT  0.0 318.32 899.4 318.88 ;
         LAYER MET3 ;
         RECT  0.0 233.68 899.4 234.24 ;
         LAYER MET3 ;
         RECT  0.0 956.8 899.4 957.36 ;
         LAYER MET3 ;
         RECT  0.0 552.0 142.24 552.56 ;
         LAYER MET4 ;
         RECT  469.2 0.0 469.76 976.68 ;
         LAYER MET4 ;
         RECT  101.2 0.0 101.76 976.68 ;
         LAYER MET3 ;
         RECT  0.0 469.2 899.4 469.76 ;
         LAYER MET3 ;
         RECT  0.0 246.56 117.4 247.12 ;
         LAYER MET3 ;
         RECT  755.32 528.08 899.4 528.64 ;
         LAYER MET3 ;
         RECT  0.0 807.76 160.64 808.32 ;
         LAYER MET3 ;
         RECT  716.68 414.0 899.4 414.56 ;
         LAYER MET4 ;
         RECT  498.64 0.0 499.2 976.68 ;
         LAYER MET3 ;
         RECT  0.0 305.44 899.4 306.0 ;
         LAYER MET4 ;
         RECT  329.36 0.0 329.92 976.68 ;
         LAYER MET4 ;
         RECT  128.8 6.44 129.36 976.68 ;
         LAYER MET4 ;
         RECT  410.32 0.0 410.88 976.68 ;
         LAYER MET3 ;
         RECT  716.68 789.36 899.4 789.92 ;
         LAYER MET3 ;
         RECT  0.0 191.36 117.4 191.92 ;
         LAYER MET4 ;
         RECT  169.28 0.0 169.84 976.68 ;
         LAYER MET4 ;
         RECT  452.64 0.0 453.2 976.68 ;
         LAYER MET3 ;
         RECT  780.16 136.16 899.4 136.72 ;
         LAYER MET3 ;
         RECT  780.16 207.92 899.4 208.48 ;
         LAYER MET3 ;
         RECT  0.0 7.36 899.4 7.92 ;
         LAYER MET4 ;
         RECT  822.48 0.0 823.04 976.68 ;
         LAYER MET3 ;
         RECT  780.16 134.32 899.4 134.88 ;
         LAYER MET3 ;
         RECT  817.88 49.68 899.4 50.24 ;
         LAYER MET3 ;
         RECT  0.0 92.0 7.0 92.56 ;
         LAYER MET3 ;
         RECT  0.0 890.56 899.4 891.12 ;
         LAYER MET3 ;
         RECT  0.0 907.12 160.64 907.68 ;
         LAYER MET4 ;
         RECT  33.12 0.0 33.68 976.68 ;
         LAYER MET3 ;
         RECT  0.0 699.2 899.4 699.76 ;
         LAYER MET4 ;
         RECT  18.4 0.0 18.96 976.68 ;
         LAYER MET3 ;
         RECT  0.0 134.32 117.4 134.88 ;
         LAYER MET4 ;
         RECT  859.28 0.0 859.84 976.68 ;
         LAYER MET3 ;
         RECT  0.0 870.32 160.64 870.88 ;
         LAYER MET4 ;
         RECT  500.48 0.0 501.04 976.68 ;
         LAYER MET3 ;
         RECT  0.0 42.32 7.0 42.88 ;
         LAYER MET4 ;
         RECT  748.88 0.0 749.44 976.68 ;
         LAYER MET3 ;
         RECT  83.72 333.04 899.4 333.6 ;
         LAYER MET3 ;
         RECT  0.0 734.16 899.4 734.72 ;
         LAYER MET4 ;
         RECT  255.76 0.0 256.32 5.16 ;
         LAYER MET3 ;
         RECT  0.0 110.4 117.4 110.96 ;
         LAYER MET4 ;
         RECT  231.84 0.0 232.4 976.68 ;
         LAYER MET3 ;
         RECT  0.0 364.32 177.2 364.88 ;
         LAYER MET3 ;
         RECT  0.0 765.44 899.4 766.0 ;
         LAYER MET3 ;
         RECT  0.0 704.72 899.4 705.28 ;
         LAYER MET4 ;
         RECT  327.52 6.44 328.08 976.68 ;
         LAYER MET3 ;
         RECT  716.68 491.28 899.4 491.84 ;
         LAYER MET3 ;
         RECT  0.0 270.48 117.4 271.04 ;
         LAYER MET3 ;
         RECT  0.0 833.52 899.4 834.08 ;
         LAYER MET3 ;
         RECT  0.0 912.64 899.4 913.2 ;
         LAYER MET3 ;
         RECT  0.0 577.76 142.24 578.32 ;
         LAYER MET4 ;
         RECT  450.8 20.24 451.36 976.68 ;
         LAYER MET4 ;
         RECT  592.48 0.0 593.04 976.68 ;
         LAYER MET4 ;
         RECT  349.6 0.0 350.16 13.44 ;
         LAYER MET4 ;
         RECT  520.72 0.0 521.28 976.68 ;
         LAYER MET3 ;
         RECT  0.0 40.48 899.4 41.04 ;
         LAYER MET4 ;
         RECT  620.08 0.0 620.64 17.12 ;
         LAYER MET3 ;
         RECT  0.0 125.12 899.4 125.68 ;
         LAYER MET4 ;
         RECT  454.48 0.0 455.04 976.68 ;
         LAYER MET3 ;
         RECT  0.0 66.24 87.96 66.8 ;
         LAYER MET4 ;
         RECT  298.08 0.0 298.64 976.68 ;
         LAYER MET4 ;
         RECT  331.2 0.0 331.76 976.68 ;
         LAYER MET3 ;
         RECT  0.0 837.2 177.2 837.76 ;
         LAYER MET3 ;
         RECT  0.0 568.56 899.4 569.12 ;
         LAYER MET4 ;
         RECT  763.6 0.0 764.16 976.68 ;
         LAYER MET4 ;
         RECT  391.92 0.0 392.48 976.68 ;
         LAYER MET4 ;
         RECT  894.24 0.0 894.8 976.68 ;
         LAYER MET3 ;
         RECT  0.0 368.0 899.4 368.56 ;
         LAYER MET3 ;
         RECT  716.68 640.32 899.4 640.88 ;
         LAYER MET3 ;
         RECT  0.0 925.52 720.0 926.08 ;
         LAYER MET4 ;
         RECT  184.0 0.0 184.56 976.68 ;
         LAYER MET4 ;
         RECT  320.16 0.0 320.72 976.68 ;
         LAYER MET4 ;
         RECT  548.32 0.0 548.88 976.68 ;
         LAYER MET3 ;
         RECT  716.68 515.2 899.4 515.76 ;
         LAYER MET3 ;
         RECT  0.0 769.12 899.4 769.68 ;
         LAYER MET3 ;
         RECT  0.0 241.04 117.4 241.6 ;
         LAYER MET4 ;
         RECT  82.8 0.0 83.36 976.68 ;
         LAYER MET4 ;
         RECT  130.64 0.0 131.2 976.68 ;
         LAYER MET3 ;
         RECT  0.0 682.64 160.64 683.2 ;
         LAYER MET3 ;
         RECT  0.0 585.12 899.4 585.68 ;
         LAYER MET3 ;
         RECT  733.24 222.64 899.4 223.2 ;
         LAYER MET3 ;
         RECT  0.0 404.8 899.4 405.36 ;
         LAYER MET3 ;
         RECT  755.32 726.8 899.4 727.36 ;
         LAYER MET3 ;
         RECT  0.0 743.36 899.4 743.92 ;
         LAYER MET3 ;
         RECT  0.0 138.0 899.4 138.56 ;
         LAYER MET3 ;
         RECT  0.0 848.24 899.4 848.8 ;
         LAYER MET4 ;
         RECT  281.52 20.24 282.08 976.68 ;
         LAYER MET4 ;
         RECT  678.96 0.0 679.52 976.68 ;
         LAYER MET4 ;
         RECT  816.96 0.0 817.52 976.68 ;
         LAYER MET3 ;
         RECT  0.0 774.64 899.4 775.2 ;
         LAYER MET3 ;
         RECT  17.48 58.88 899.4 59.44 ;
         LAYER MET3 ;
         RECT  0.0 929.2 899.4 929.76 ;
         LAYER MET3 ;
         RECT  0.0 379.04 142.24 379.6 ;
         LAYER MET4 ;
         RECT  106.72 0.0 107.28 976.68 ;
         LAYER MET3 ;
         RECT  0.0 299.92 80.6 300.48 ;
         LAYER MET4 ;
         RECT  513.36 0.0 513.92 976.68 ;
         LAYER MET3 ;
         RECT  716.68 638.48 899.4 639.04 ;
         LAYER MET3 ;
         RECT  731.4 408.48 899.4 409.04 ;
         LAYER MET4 ;
         RECT  384.56 0.0 385.12 976.68 ;
         LAYER MET3 ;
         RECT  0.0 349.6 899.4 350.16 ;
         LAYER MET3 ;
         RECT  0.0 331.2 899.4 331.76 ;
         LAYER MET4 ;
         RECT  881.36 0.0 881.92 976.68 ;
         LAYER MET4 ;
         RECT  301.76 0.0 302.32 976.68 ;
         LAYER MET4 ;
         RECT  802.24 0.0 802.8 976.68 ;
         LAYER MET3 ;
         RECT  0.0 544.64 899.4 545.2 ;
         LAYER MET3 ;
         RECT  0.0 345.92 899.4 346.48 ;
         LAYER MET4 ;
         RECT  818.8 64.4 819.36 976.68 ;
         LAYER MET4 ;
         RECT  160.08 6.44 160.64 976.68 ;
         LAYER MET4 ;
         RECT  226.32 6.44 226.88 976.68 ;
         LAYER MET4 ;
         RECT  690.0 0.0 690.56 976.68 ;
         LAYER MET3 ;
         RECT  0.0 712.08 899.4 712.64 ;
         LAYER MET3 ;
         RECT  733.24 794.88 899.4 795.44 ;
         LAYER MET3 ;
         RECT  0.0 546.48 160.64 547.04 ;
         LAYER MET3 ;
         RECT  0.0 561.2 899.4 561.76 ;
         LAYER MET4 ;
         RECT  445.28 0.0 445.84 976.68 ;
         LAYER MET3 ;
         RECT  0.0 51.52 28.16 52.08 ;
         LAYER MET3 ;
         RECT  0.0 106.72 117.4 107.28 ;
         LAYER MET4 ;
         RECT  669.76 0.0 670.32 976.68 ;
         LAYER MET4 ;
         RECT  235.52 0.0 236.08 976.68 ;
         LAYER MET3 ;
         RECT  0.0 397.44 160.64 398.0 ;
         LAYER MET4 ;
         RECT  77.28 0.0 77.84 976.68 ;
         LAYER MET3 ;
         RECT  0.0 237.36 899.4 237.92 ;
         LAYER MET3 ;
         RECT  716.68 217.12 899.4 217.68 ;
         LAYER MET3 ;
         RECT  0.0 29.44 899.4 30.0 ;
         LAYER MET3 ;
         RECT  0.0 715.76 899.4 716.32 ;
         LAYER MET4 ;
         RECT  721.28 0.0 721.84 976.68 ;
         LAYER MET3 ;
         RECT  716.68 787.52 899.4 788.08 ;
         LAYER MET3 ;
         RECT  0.0 763.6 177.2 764.16 ;
         LAYER MET4 ;
         RECT  255.76 12.88 256.32 976.68 ;
         LAYER MET4 ;
         RECT  272.32 0.0 272.88 5.16 ;
         LAYER MET3 ;
         RECT  405.72 5.52 899.4 6.08 ;
         LAYER MET3 ;
         RECT  716.68 539.12 899.4 539.68 ;
         LAYER MET3 ;
         RECT  716.68 588.8 899.4 589.36 ;
         LAYER MET4 ;
         RECT  620.08 20.24 620.64 976.68 ;
         LAYER MET4 ;
         RECT  489.44 0.0 490.0 976.68 ;
         LAYER MET3 ;
         RECT  810.52 938.4 899.4 938.96 ;
         LAYER MET4 ;
         RECT  697.36 0.0 697.92 976.68 ;
         LAYER MET3 ;
         RECT  716.68 737.84 899.4 738.4 ;
         LAYER MET4 ;
         RECT  108.56 0.0 109.12 976.68 ;
         LAYER MET3 ;
         RECT  0.0 550.16 899.4 550.72 ;
         LAYER MET3 ;
         RECT  0.0 500.48 899.4 501.04 ;
         LAYER MET3 ;
         RECT  0.0 230.0 899.4 230.56 ;
         LAYER MET3 ;
         RECT  0.0 658.72 160.64 659.28 ;
         LAYER MET3 ;
         RECT  755.32 750.72 899.4 751.28 ;
         LAYER MET4 ;
         RECT  44.16 0.0 44.72 976.68 ;
         LAYER MET4 ;
         RECT  610.88 0.0 611.44 976.68 ;
         LAYER MET4 ;
         RECT  68.08 0.0 68.64 976.68 ;
         LAYER MET3 ;
         RECT  0.0 966.0 749.44 966.56 ;
         LAYER MET4 ;
         RECT  734.16 0.0 734.72 976.68 ;
         LAYER MET4 ;
         RECT  99.36 0.0 99.92 976.68 ;
         LAYER MET3 ;
         RECT  0.0 22.08 179.04 22.64 ;
         LAYER MET3 ;
         RECT  0.0 132.48 117.4 133.04 ;
         LAYER MET3 ;
         RECT  780.16 185.84 899.4 186.4 ;
         LAYER MET3 ;
         RECT  0.0 800.4 142.24 800.96 ;
         LAYER MET4 ;
         RECT  609.04 0.0 609.6 976.68 ;
         LAYER MET3 ;
         RECT  0.0 747.04 899.4 747.6 ;
         LAYER MET3 ;
         RECT  0.0 218.96 899.4 219.52 ;
         LAYER MET4 ;
         RECT  152.72 0.0 153.28 976.68 ;
         LAYER MET3 ;
         RECT  0.0 796.72 899.4 797.28 ;
         LAYER MET3 ;
         RECT  0.0 158.24 899.4 158.8 ;
         LAYER MET3 ;
         RECT  0.0 408.48 162.48 409.04 ;
         LAYER MET4 ;
         RECT  671.6 0.0 672.16 976.68 ;
         LAYER MET4 ;
         RECT  172.96 0.0 173.52 5.16 ;
         LAYER MET3 ;
         RECT  0.0 226.32 899.4 226.88 ;
         LAYER MET3 ;
         RECT  0.0 235.52 160.64 236.08 ;
         LAYER MET4 ;
         RECT  752.56 0.0 753.12 976.68 ;
         LAYER MET3 ;
         RECT  0.0 736.0 899.4 736.56 ;
         LAYER MET4 ;
         RECT  644.0 0.0 644.56 976.68 ;
         LAYER MET4 ;
         RECT  787.52 0.0 788.08 976.68 ;
         LAYER MET3 ;
         RECT  716.68 314.64 899.4 315.2 ;
         LAYER MET4 ;
         RECT  126.96 0.0 127.52 976.68 ;
         LAYER MET4 ;
         RECT  877.68 0.0 878.24 976.68 ;
         LAYER MET4 ;
         RECT  371.68 18.4 372.24 976.68 ;
         LAYER MET3 ;
         RECT  780.16 206.08 899.4 206.64 ;
         LAYER MET3 ;
         RECT  874.0 962.32 899.4 962.88 ;
         LAYER MET4 ;
         RECT  588.8 0.0 589.36 976.68 ;
         LAYER MET4 ;
         RECT  839.04 0.0 839.6 976.68 ;
         LAYER MET4 ;
         RECT  119.6 0.0 120.16 976.68 ;
         LAYER MET3 ;
         RECT  0.0 614.56 899.4 615.12 ;
         LAYER MET4 ;
         RECT  239.2 14.72 239.76 976.68 ;
         LAYER MET4 ;
         RECT  474.72 0.0 475.28 976.68 ;
         LAYER MET4 ;
         RECT  287.04 0.0 287.6 976.68 ;
         LAYER MET3 ;
         RECT  0.0 426.88 899.4 427.44 ;
         LAYER MET4 ;
         RECT  156.4 0.0 156.96 5.16 ;
         LAYER MET3 ;
         RECT  780.16 257.6 899.4 258.16 ;
         LAYER MET3 ;
         RECT  780.16 268.64 899.4 269.2 ;
         LAYER MET4 ;
         RECT  246.56 0.0 247.12 9.76 ;
         LAYER MET4 ;
         RECT  200.56 0.0 201.12 976.68 ;
         LAYER MET4 ;
         RECT  401.12 0.0 401.68 976.68 ;
         LAYER MET3 ;
         RECT  716.68 690.0 899.4 690.56 ;
         LAYER MET3 ;
         RECT  0.0 123.28 117.4 123.84 ;
         LAYER MET3 ;
         RECT  0.0 529.92 899.4 530.48 ;
         LAYER MET4 ;
         RECT  189.52 0.0 190.08 5.16 ;
         LAYER MET3 ;
         RECT  0.0 322.0 160.64 322.56 ;
         LAYER MET3 ;
         RECT  91.08 66.24 899.4 66.8 ;
         LAYER MET4 ;
         RECT  695.52 0.0 696.08 976.68 ;
         LAYER MET3 ;
         RECT  733.24 596.16 899.4 596.72 ;
         LAYER MET3 ;
         RECT  19.32 103.04 899.4 103.6 ;
         LAYER MET3 ;
         RECT  0.0 320.16 77.84 320.72 ;
         LAYER MET3 ;
         RECT  0.0 805.92 899.4 806.48 ;
         LAYER MET4 ;
         RECT  9.2 0.0 9.76 976.68 ;
         LAYER MET4 ;
         RECT  14.72 0.0 15.28 976.68 ;
         LAYER MET4 ;
         RECT  92.0 0.0 92.56 976.68 ;
         LAYER MET3 ;
         RECT  733.24 149.04 899.4 149.6 ;
         LAYER MET3 ;
         RECT  0.0 618.24 899.4 618.8 ;
         LAYER MET4 ;
         RECT  3.68 0.0 4.24 976.68 ;
         LAYER MET3 ;
         RECT  0.0 791.2 899.4 791.76 ;
         LAYER MET3 ;
         RECT  0.0 892.4 753.12 892.96 ;
         LAYER MET3 ;
         RECT  0.0 147.2 899.4 147.76 ;
         LAYER MET3 ;
         RECT  0.0 476.56 899.4 477.12 ;
         LAYER MET4 ;
         RECT  793.04 0.0 793.6 976.68 ;
         LAYER MET3 ;
         RECT  733.24 857.44 899.4 858.0 ;
         LAYER MET3 ;
         RECT  0.0 231.84 899.4 232.4 ;
         LAYER MET4 ;
         RECT  344.08 6.44 344.64 976.68 ;
         LAYER MET3 ;
         RECT  0.0 340.4 177.2 340.96 ;
         LAYER MET3 ;
         RECT  0.0 33.12 87.96 33.68 ;
         LAYER MET3 ;
         RECT  0.0 90.16 806.48 90.72 ;
         LAYER MET4 ;
         RECT  518.88 20.24 519.44 976.68 ;
         LAYER MET3 ;
         RECT  0.0 509.68 162.48 510.24 ;
         LAYER MET4 ;
         RECT  511.52 0.0 512.08 976.68 ;
         LAYER MET3 ;
         RECT  733.24 658.72 899.4 659.28 ;
         LAYER MET3 ;
         RECT  716.68 713.92 899.4 714.48 ;
         LAYER MET3 ;
         RECT  0.0 402.96 142.24 403.52 ;
         LAYER MET3 ;
         RECT  0.0 434.24 160.64 434.8 ;
         LAYER MET3 ;
         RECT  716.68 864.8 899.4 865.36 ;
         LAYER MET4 ;
         RECT  844.56 0.0 845.12 976.68 ;
         LAYER MET4 ;
         RECT  259.44 0.0 260.0 976.68 ;
         LAYER MET4 ;
         RECT  570.4 0.0 570.96 976.68 ;
         LAYER MET4 ;
         RECT  103.04 0.0 103.6 976.68 ;
         LAYER MET4 ;
         RECT  625.6 0.0 626.16 976.68 ;
         LAYER MET3 ;
         RECT  0.0 517.04 899.4 517.6 ;
         LAYER MET3 ;
         RECT  892.4 897.92 899.4 898.48 ;
         LAYER MET4 ;
         RECT  279.68 0.0 280.24 962.88 ;
         LAYER MET4 ;
         RECT  288.88 14.72 289.44 976.68 ;
         LAYER MET3 ;
         RECT  0.0 34.96 899.4 35.52 ;
         LAYER MET3 ;
         RECT  0.0 840.88 899.4 841.44 ;
         LAYER MET3 ;
         RECT  723.12 916.32 899.4 916.88 ;
         LAYER MET3 ;
         RECT  0.0 780.16 899.4 780.72 ;
         LAYER MET4 ;
         RECT  583.28 0.0 583.84 976.68 ;
         LAYER MET3 ;
         RECT  0.0 287.04 899.4 287.6 ;
         LAYER MET3 ;
         RECT  0.0 518.88 899.4 519.44 ;
         LAYER MET3 ;
         RECT  892.4 881.36 899.4 881.92 ;
         LAYER MET3 ;
         RECT  0.0 425.04 899.4 425.6 ;
         LAYER MET4 ;
         RECT  386.4 0.0 386.96 976.68 ;
         LAYER MET4 ;
         RECT  765.44 0.0 766.0 976.68 ;
         LAYER MET3 ;
         RECT  0.0 866.64 899.4 867.2 ;
         LAYER MET4 ;
         RECT  789.36 0.0 789.92 976.68 ;
         LAYER MET4 ;
         RECT  713.92 0.0 714.48 976.68 ;
         LAYER MET3 ;
         RECT  0.0 590.64 177.2 591.2 ;
         LAYER MET3 ;
         RECT  0.0 596.16 160.64 596.72 ;
         LAYER MET4 ;
         RECT  888.72 0.0 889.28 976.68 ;
         LAYER MET3 ;
         RECT  733.24 235.52 899.4 236.08 ;
         LAYER MET4 ;
         RECT  875.84 0.0 876.4 976.68 ;
         LAYER MET3 ;
         RECT  0.0 793.04 899.4 793.6 ;
         LAYER MET4 ;
         RECT  809.6 0.0 810.16 976.68 ;
         LAYER MET3 ;
         RECT  0.0 472.88 899.4 473.44 ;
         LAYER MET4 ;
         RECT  732.32 0.0 732.88 976.68 ;
         LAYER MET4 ;
         RECT  835.36 0.0 835.92 976.68 ;
         LAYER MET4 ;
         RECT  857.44 0.0 858.0 976.68 ;
         LAYER MET4 ;
         RECT  196.88 0.0 197.44 976.68 ;
         LAYER MET4 ;
         RECT  826.16 0.0 826.72 976.68 ;
         LAYER MET3 ;
         RECT  0.0 975.2 899.4 975.76 ;
         LAYER MET4 ;
         RECT  233.68 0.0 234.24 976.68 ;
         LAYER MET3 ;
         RECT  0.0 642.16 899.4 642.72 ;
         LAYER MET4 ;
         RECT  377.2 6.44 377.76 976.68 ;
         LAYER MET3 ;
         RECT  0.0 119.6 117.4 120.16 ;
         LAYER MET4 ;
         RECT  220.8 0.0 221.36 976.68 ;
         LAYER MET4 ;
         RECT  846.4 0.0 846.96 976.68 ;
         LAYER MET4 ;
         RECT  533.6 0.0 534.16 976.68 ;
         LAYER MET4 ;
         RECT  649.52 0.0 650.08 976.68 ;
         LAYER MET3 ;
         RECT  0.0 145.36 899.4 145.92 ;
         LAYER MET4 ;
         RECT  338.56 0.0 339.12 5.16 ;
         LAYER MET3 ;
         RECT  0.0 285.2 117.4 285.76 ;
         LAYER MET3 ;
         RECT  0.0 471.04 160.64 471.6 ;
         LAYER MET4 ;
         RECT  575.92 0.0 576.48 976.68 ;
         LAYER MET4 ;
         RECT  230.0 0.0 230.56 976.68 ;
         LAYER MET3 ;
         RECT  0.0 428.72 142.24 429.28 ;
         LAYER MET3 ;
         RECT  0.0 117.76 117.4 118.32 ;
         LAYER MET3 ;
         RECT  733.24 371.68 899.4 372.24 ;
         LAYER MET4 ;
         RECT  853.76 0.0 854.32 976.68 ;
         LAYER MET4 ;
         RECT  360.64 6.44 361.2 976.68 ;
         LAYER MET4 ;
         RECT  395.6 0.0 396.16 976.68 ;
         LAYER MET3 ;
         RECT  0.0 360.64 899.4 361.2 ;
         LAYER MET3 ;
         RECT  0.0 375.36 899.4 375.92 ;
         LAYER MET4 ;
         RECT  636.64 0.0 637.2 976.68 ;
         LAYER MET3 ;
         RECT  0.0 272.32 117.4 272.88 ;
         LAYER MET4 ;
         RECT  813.28 0.0 813.84 976.68 ;
         LAYER MET3 ;
         RECT  0.0 673.44 899.4 674.0 ;
         LAYER MET3 ;
         RECT  43.24 20.24 899.4 20.8 ;
         LAYER MET3 ;
         RECT  0.0 667.92 899.4 668.48 ;
         LAYER MET3 ;
         RECT  780.16 193.2 899.4 193.76 ;
         LAYER MET4 ;
         RECT  596.16 0.0 596.72 976.68 ;
         LAYER MET4 ;
         RECT  850.08 0.0 850.64 976.68 ;
         LAYER MET3 ;
         RECT  733.24 334.88 899.4 335.44 ;
         LAYER MET4 ;
         RECT  872.16 0.0 872.72 976.68 ;
         LAYER MET3 ;
         RECT  780.16 121.44 899.4 122.0 ;
         LAYER MET3 ;
         RECT  0.0 524.4 899.4 524.96 ;
         LAYER MET3 ;
         RECT  0.0 632.96 160.64 633.52 ;
         LAYER MET4 ;
         RECT  417.68 0.0 418.24 976.68 ;
         LAYER MET4 ;
         RECT  883.2 0.0 883.76 976.68 ;
         LAYER MET3 ;
         RECT  0.0 684.48 899.4 685.04 ;
         LAYER MET4 ;
         RECT  824.32 0.0 824.88 976.68 ;
         LAYER MET3 ;
         RECT  780.16 195.04 899.4 195.6 ;
         LAYER MET4 ;
         RECT  42.32 0.0 42.88 976.68 ;
         LAYER MET4 ;
         RECT  441.6 0.0 442.16 976.68 ;
         LAYER MET3 ;
         RECT  755.32 478.4 899.4 478.96 ;
         LAYER MET4 ;
         RECT  737.84 0.0 738.4 976.68 ;
         LAYER MET4 ;
         RECT  217.12 0.0 217.68 976.68 ;
         LAYER MET3 ;
         RECT  733.24 483.92 899.4 484.48 ;
         LAYER MET4 ;
         RECT  202.4 0.0 202.96 976.68 ;
         LAYER MET3 ;
         RECT  0.0 528.08 142.24 528.64 ;
         LAYER MET4 ;
         RECT  57.04 0.0 57.6 976.68 ;
         LAYER MET3 ;
         RECT  0.0 625.6 899.4 626.16 ;
         LAYER MET4 ;
         RECT  209.76 6.44 210.32 976.68 ;
         LAYER MET4 ;
         RECT  423.2 0.0 423.76 976.68 ;
         LAYER MET3 ;
         RECT  0.0 857.44 160.64 858.0 ;
         LAYER MET3 ;
         RECT  0.0 616.4 899.4 616.96 ;
         LAYER MET3 ;
         RECT  0.0 564.88 899.4 565.44 ;
         LAYER MET3 ;
         RECT  0.0 923.68 899.4 924.24 ;
         LAYER MET4 ;
         RECT  139.84 0.0 140.4 976.68 ;
         LAYER MET3 ;
         RECT  0.0 215.28 177.2 215.84 ;
         LAYER MET3 ;
         RECT  0.0 3.68 89.8 4.24 ;
         LAYER MET4 ;
         RECT  318.32 0.0 318.88 976.68 ;
         LAYER MET3 ;
         RECT  780.16 119.6 899.4 120.16 ;
         LAYER MET3 ;
         RECT  0.0 454.48 899.4 455.04 ;
         LAYER MET3 ;
         RECT  0.0 649.52 899.4 650.08 ;
         LAYER MET3 ;
         RECT  716.68 688.16 899.4 688.72 ;
         LAYER MET4 ;
         RECT  147.2 0.0 147.76 976.68 ;
         LAYER MET3 ;
         RECT  733.24 645.84 899.4 646.4 ;
         LAYER MET3 ;
         RECT  0.0 680.8 899.4 681.36 ;
         LAYER MET4 ;
         RECT  1.84 114.08 2.4 976.68 ;
         LAYER MET4 ;
         RECT  5.52 0.0 6.08 976.68 ;
         LAYER MET3 ;
         RECT  780.16 130.64 899.4 131.2 ;
         LAYER MET3 ;
         RECT  0.0 452.64 142.24 453.2 ;
         LAYER MET4 ;
         RECT  428.72 0.0 429.28 976.68 ;
         LAYER MET4 ;
         RECT  688.16 20.24 688.72 976.68 ;
         LAYER MET3 ;
         RECT  716.68 590.64 899.4 591.2 ;
         LAYER MET3 ;
         RECT  0.0 185.84 117.4 186.4 ;
         LAYER MET4 ;
         RECT  268.64 0.0 269.2 976.68 ;
         LAYER MET3 ;
         RECT  755.32 154.56 899.4 155.12 ;
         LAYER MET3 ;
         RECT  0.0 450.8 899.4 451.36 ;
         LAYER MET4 ;
         RECT  222.64 12.88 223.2 976.68 ;
         LAYER MET4 ;
         RECT  185.84 0.0 186.4 976.68 ;
         LAYER MET3 ;
         RECT  0.0 255.76 117.4 256.32 ;
         LAYER MET4 ;
         RECT  264.96 0.0 265.52 976.68 ;
         LAYER MET3 ;
         RECT  0.0 224.48 899.4 225.04 ;
         LAYER MET3 ;
         RECT  733.24 298.08 899.4 298.64 ;
         LAYER MET3 ;
         RECT  733.24 782.0 899.4 782.56 ;
         LAYER MET3 ;
         RECT  0.0 809.6 899.4 810.16 ;
         LAYER MET3 ;
         RECT  809.6 934.72 899.4 935.28 ;
         LAYER MET3 ;
         RECT  0.0 967.84 899.4 968.4 ;
         LAYER MET4 ;
         RECT  64.4 0.0 64.96 976.68 ;
         LAYER MET3 ;
         RECT  808.68 973.36 899.4 973.92 ;
         LAYER MET3 ;
         RECT  716.68 316.48 899.4 317.04 ;
         LAYER MET3 ;
         RECT  0.0 702.88 899.4 703.44 ;
         LAYER MET3 ;
         RECT  733.24 546.48 899.4 547.04 ;
         LAYER MET4 ;
         RECT  805.92 0.0 806.48 976.68 ;
         LAYER MET3 ;
         RECT  0.0 23.92 899.4 24.48 ;
         LAYER MET3 ;
         RECT  0.0 621.92 899.4 622.48 ;
         LAYER MET3 ;
         RECT  0.0 38.64 89.8 39.2 ;
         LAYER MET3 ;
         RECT  733.24 732.32 899.4 732.88 ;
         LAYER MET4 ;
         RECT  193.2 0.0 193.76 976.68 ;
         LAYER MET3 ;
         RECT  0.0 723.12 899.4 723.68 ;
         LAYER MET3 ;
         RECT  716.68 141.68 899.4 142.24 ;
         LAYER MET3 ;
         RECT  733.24 844.56 899.4 845.12 ;
         LAYER MET3 ;
         RECT  780.16 283.36 899.4 283.92 ;
         LAYER MET3 ;
         RECT  0.0 557.52 899.4 558.08 ;
         LAYER MET4 ;
         RECT  36.8 12.88 37.36 976.68 ;
         LAYER MET4 ;
         RECT  174.8 0.0 175.36 976.68 ;
         LAYER MET4 ;
         RECT  393.76 6.44 394.32 976.68 ;
         LAYER MET3 ;
         RECT  0.0 298.08 160.64 298.64 ;
         LAYER MET3 ;
         RECT  0.0 99.36 160.64 99.92 ;
         LAYER MET4 ;
         RECT  388.24 0.0 388.8 5.16 ;
         LAYER MET3 ;
         RECT  0.0 406.64 899.4 407.2 ;
         LAYER MET3 ;
         RECT  0.0 419.52 899.4 420.08 ;
         LAYER MET3 ;
         RECT  0.0 198.72 160.64 199.28 ;
         LAYER MET4 ;
         RECT  79.12 0.0 79.68 976.68 ;
         LAYER MET3 ;
         RECT  0.0 824.32 899.4 824.88 ;
         LAYER MET3 ;
         RECT  0.0 563.04 899.4 563.6 ;
         LAYER MET4 ;
         RECT  717.6 0.0 718.16 976.68 ;
         LAYER MET3 ;
         RECT  0.0 384.56 160.64 385.12 ;
         LAYER MET3 ;
         RECT  755.32 303.6 899.4 304.16 ;
         LAYER MET3 ;
         RECT  0.0 489.44 177.2 490.0 ;
         LAYER MET3 ;
         RECT  733.24 570.4 899.4 570.96 ;
         LAYER MET4 ;
         RECT  660.56 0.0 661.12 976.68 ;
         LAYER MET4 ;
         RECT  623.76 0.0 624.32 976.68 ;
         LAYER MET3 ;
         RECT  817.88 68.08 899.4 68.64 ;
         LAYER MET3 ;
         RECT  0.0 883.2 899.4 883.76 ;
         LAYER MET4 ;
         RECT  885.04 0.0 885.6 976.68 ;
         LAYER MET3 ;
         RECT  0.0 75.44 7.0 76.0 ;
         LAYER MET3 ;
         RECT  0.0 432.4 899.4 432.96 ;
         LAYER MET3 ;
         RECT  733.24 99.36 899.4 99.92 ;
         LAYER MET3 ;
         RECT  0.0 366.16 177.2 366.72 ;
         LAYER MET3 ;
         RECT  0.0 605.36 899.4 605.92 ;
         LAYER MET3 ;
         RECT  755.32 552.0 899.4 552.56 ;
         LAYER MET3 ;
         RECT  451.72 12.88 899.4 13.44 ;
         LAYER MET4 ;
         RECT  66.24 0.0 66.8 976.68 ;
         LAYER MET3 ;
         RECT  0.0 485.76 899.4 486.32 ;
         LAYER MET4 ;
         RECT  222.64 0.0 223.2 5.16 ;
         LAYER MET4 ;
         RECT  675.28 0.0 675.84 976.68 ;
         LAYER MET4 ;
         RECT  456.32 0.0 456.88 976.68 ;
         LAYER MET3 ;
         RECT  0.0 47.84 121.08 48.4 ;
         LAYER MET3 ;
         RECT  0.0 377.2 899.4 377.76 ;
         LAYER MET3 ;
         RECT  797.64 253.92 899.4 254.48 ;
         LAYER MET3 ;
         RECT  132.48 47.84 899.4 48.4 ;
         LAYER MET3 ;
         RECT  0.0 598.0 899.4 598.56 ;
         LAYER MET4 ;
         RECT  34.96 0.0 35.52 976.68 ;
         LAYER MET3 ;
         RECT  0.0 283.36 117.4 283.92 ;
         LAYER MET3 ;
         RECT  780.16 172.96 899.4 173.52 ;
         LAYER MET3 ;
         RECT  0.0 312.8 88.88 313.36 ;
         LAYER MET3 ;
         RECT  0.0 566.72 899.4 567.28 ;
         LAYER MET4 ;
         RECT  7.36 0.0 7.92 976.68 ;
         LAYER MET3 ;
         RECT  0.0 445.28 899.4 445.84 ;
         LAYER MET4 ;
         RECT  439.76 0.0 440.32 976.68 ;
         LAYER MET3 ;
         RECT  0.0 204.24 100.84 204.8 ;
         LAYER MET4 ;
         RECT  114.08 0.0 114.64 976.68 ;
         LAYER MET3 ;
         RECT  0.0 207.92 117.4 208.48 ;
         LAYER MET3 ;
         RECT  797.64 178.48 899.4 179.04 ;
         LAYER MET3 ;
         RECT  0.0 156.4 899.4 156.96 ;
         LAYER MET3 ;
         RECT  0.0 520.72 160.64 521.28 ;
         LAYER MET3 ;
         RECT  0.0 391.92 177.2 392.48 ;
         LAYER MET3 ;
         RECT  0.0 570.4 160.64 570.96 ;
         LAYER MET3 ;
         RECT  716.68 763.6 899.4 764.16 ;
         LAYER MET4 ;
         RECT  104.88 0.0 105.44 976.68 ;
         LAYER MET3 ;
         RECT  98.44 336.72 899.4 337.28 ;
         LAYER MET4 ;
         RECT  691.84 0.0 692.4 976.68 ;
         LAYER MET4 ;
         RECT  673.44 0.0 674.0 976.68 ;
         LAYER MET3 ;
         RECT  810.52 921.84 899.4 922.4 ;
         LAYER MET3 ;
         RECT  0.0 141.68 177.2 142.24 ;
         LAYER MET3 ;
         RECT  731.4 770.96 899.4 771.52 ;
         LAYER MET4 ;
         RECT  355.12 14.72 355.68 976.68 ;
         LAYER MET4 ;
         RECT  831.68 0.0 832.24 976.68 ;
         LAYER MET4 ;
         RECT  704.72 0.0 705.28 976.68 ;
         LAYER MET3 ;
         RECT  0.0 290.72 177.2 291.28 ;
         LAYER MET3 ;
         RECT  755.32 452.64 899.4 453.2 ;
         LAYER MET4 ;
         RECT  195.04 6.44 195.6 976.68 ;
         LAYER MET4 ;
         RECT  577.76 0.0 578.32 976.68 ;
         LAYER MET4 ;
         RECT  274.16 0.0 274.72 976.68 ;
         LAYER MET4 ;
         RECT  627.44 0.0 628.0 976.68 ;
         LAYER MET4 ;
         RECT  502.32 0.0 502.88 976.68 ;
         LAYER MET4 ;
         RECT  528.08 0.0 528.64 976.68 ;
         LAYER MET3 ;
         RECT  0.0 220.8 899.4 221.36 ;
         LAYER MET4 ;
         RECT  759.92 0.0 760.48 976.68 ;
         LAYER MET4 ;
         RECT  686.32 0.0 686.88 962.88 ;
         LAYER MET4 ;
         RECT  88.32 0.0 88.88 976.68 ;
         LAYER MET3 ;
         RECT  0.0 436.08 899.4 436.64 ;
         LAYER MET3 ;
         RECT  0.0 675.28 899.4 675.84 ;
         LAYER MET3 ;
         RECT  755.32 701.04 899.4 701.6 ;
         LAYER MET3 ;
         RECT  755.32 899.76 899.4 900.32 ;
         LAYER MET3 ;
         RECT  552.92 16.56 899.4 17.12 ;
         LAYER MET4 ;
         RECT  69.92 0.0 70.48 976.68 ;
         LAYER MET3 ;
         RECT  0.0 180.32 117.4 180.88 ;
         LAYER MET4 ;
         RECT  616.4 0.0 616.96 962.88 ;
         LAYER MET4 ;
         RECT  261.28 6.44 261.84 976.68 ;
         LAYER MET3 ;
         RECT  780.16 171.12 899.4 171.68 ;
         LAYER MET3 ;
         RECT  0.0 211.6 899.4 212.16 ;
         LAYER MET4 ;
         RECT  461.84 0.0 462.4 976.68 ;
         LAYER MET4 ;
         RECT  614.56 0.0 615.12 976.68 ;
         LAYER MET3 ;
         RECT  0.0 31.28 121.08 31.84 ;
         LAYER MET4 ;
         RECT  53.36 0.0 53.92 976.68 ;
         LAYER MET4 ;
         RECT  581.44 0.0 582.0 976.68 ;
         LAYER MET3 ;
         RECT  0.0 467.36 899.4 467.92 ;
         LAYER MET3 ;
         RECT  0.0 502.32 142.24 502.88 ;
         LAYER MET3 ;
         RECT  733.24 695.52 899.4 696.08 ;
         LAYER MET3 ;
         RECT  0.0 713.92 177.2 714.48 ;
         LAYER MET3 ;
         RECT  0.0 388.24 899.4 388.8 ;
         LAYER MET3 ;
         RECT  0.0 439.76 177.2 440.32 ;
         LAYER MET4 ;
         RECT  242.88 0.0 243.44 976.68 ;
         LAYER MET4 ;
         RECT  774.64 0.0 775.2 976.68 ;
         LAYER MET3 ;
         RECT  755.32 577.76 899.4 578.32 ;
         LAYER MET3 ;
         RECT  0.0 846.4 899.4 846.96 ;
         LAYER MET4 ;
         RECT  770.96 0.0 771.52 970.24 ;
         LAYER MET3 ;
         RECT  733.24 496.8 899.4 497.36 ;
         LAYER MET3 ;
         RECT  755.32 850.08 899.4 850.64 ;
         LAYER MET4 ;
         RECT  656.88 0.0 657.44 976.68 ;
         LAYER MET3 ;
         RECT  0.0 610.88 899.4 611.44 ;
         LAYER MET3 ;
         RECT  716.68 264.96 899.4 265.52 ;
         LAYER MET3 ;
         RECT  780.16 117.76 899.4 118.32 ;
         LAYER MET3 ;
         RECT  0.0 417.68 899.4 418.24 ;
         LAYER MET4 ;
         RECT  590.64 0.0 591.2 976.68 ;
         LAYER MET4 ;
         RECT  897.92 926.44 898.48 976.68 ;
         LAYER MET3 ;
         RECT  0.0 931.04 882.84 931.6 ;
         LAYER MET3 ;
         RECT  0.0 506.0 899.4 506.56 ;
         LAYER MET3 ;
         RECT  0.0 874.0 899.4 874.56 ;
         LAYER MET3 ;
         RECT  780.16 241.04 899.4 241.6 ;
         LAYER MET3 ;
         RECT  733.24 347.76 899.4 348.32 ;
         LAYER MET3 ;
         RECT  0.0 908.96 881.0 909.52 ;
         LAYER MET4 ;
         RECT  167.44 0.0 168.0 976.68 ;
         LAYER MET4 ;
         RECT  471.04 0.0 471.6 976.68 ;
         LAYER MET4 ;
         RECT  561.2 0.0 561.76 976.68 ;
         LAYER MET3 ;
         RECT  0.0 875.84 142.24 876.4 ;
         LAYER MET4 ;
         RECT  796.72 0.0 797.28 976.68 ;
         LAYER MET3 ;
         RECT  0.0 942.08 899.4 942.64 ;
         LAYER MET3 ;
         RECT  0.0 631.12 899.4 631.68 ;
         LAYER MET4 ;
         RECT  436.08 0.0 436.64 976.68 ;
         LAYER MET3 ;
         RECT  0.0 818.8 899.4 819.36 ;
         LAYER MET4 ;
         RECT  294.4 6.44 294.96 976.68 ;
         LAYER MET3 ;
         RECT  0.0 248.4 160.64 248.96 ;
         LAYER MET3 ;
         RECT  0.0 686.32 899.4 686.88 ;
         LAYER MET3 ;
         RECT  771.88 971.52 899.4 972.08 ;
         LAYER MET3 ;
         RECT  780.16 182.16 899.4 182.72 ;
         LAYER MET3 ;
         RECT  755.32 379.04 899.4 379.6 ;
         LAYER MET3 ;
         RECT  0.0 97.52 117.4 98.08 ;
         LAYER MET4 ;
         RECT  463.68 0.0 464.24 976.68 ;
         LAYER MET3 ;
         RECT  0.0 463.68 899.4 464.24 ;
         LAYER MET3 ;
         RECT  0.0 888.72 177.2 889.28 ;
         LAYER MET4 ;
         RECT  566.72 0.0 567.28 976.68 ;
         LAYER MET3 ;
         RECT  0.0 901.6 881.0 902.16 ;
         LAYER MET3 ;
         RECT  0.0 586.96 899.4 587.52 ;
         LAYER MET4 ;
         RECT  206.08 0.0 206.64 5.16 ;
         LAYER MET3 ;
         RECT  716.68 415.84 899.4 416.4 ;
         LAYER MET3 ;
         RECT  0.0 77.28 899.4 77.84 ;
         LAYER MET3 ;
         RECT  716.68 366.16 899.4 366.72 ;
         LAYER MET3 ;
         RECT  0.0 660.56 899.4 661.12 ;
         LAYER MET4 ;
         RECT  568.56 0.0 569.12 976.68 ;
         LAYER MET4 ;
         RECT  829.84 0.0 830.4 976.68 ;
         LAYER MET3 ;
         RECT  0.0 25.76 899.4 26.32 ;
         LAYER MET4 ;
         RECT  870.32 0.0 870.88 976.68 ;
         LAYER MET3 ;
         RECT  0.0 344.08 899.4 344.64 ;
         LAYER MET3 ;
         RECT  0.0 130.64 117.4 131.2 ;
         LAYER MET3 ;
         RECT  0.0 962.32 176.28 962.88 ;
         LAYER MET4 ;
         RECT  458.16 0.0 458.72 976.68 ;
         LAYER MET3 ;
         RECT  716.68 837.2 899.4 837.76 ;
         LAYER MET4 ;
         RECT  244.72 6.44 245.28 976.68 ;
         LAYER MET4 ;
         RECT  552.0 0.0 552.56 15.28 ;
         LAYER MET3 ;
         RECT  0.0 393.76 899.4 394.32 ;
         LAYER MET4 ;
         RECT  266.8 0.0 267.36 976.68 ;
         LAYER MET3 ;
         RECT  0.0 539.12 177.2 539.68 ;
         LAYER MET4 ;
         RECT  658.72 0.0 659.28 976.68 ;
         LAYER MET3 ;
         RECT  0.0 656.88 899.4 657.44 ;
         LAYER MET3 ;
         RECT  0.0 905.28 899.4 905.84 ;
         LAYER MET3 ;
         RECT  19.32 112.24 899.4 112.8 ;
         LAYER MET3 ;
         RECT  716.68 441.6 899.4 442.16 ;
         LAYER MET3 ;
         RECT  0.0 296.24 899.4 296.8 ;
         LAYER MET4 ;
         RECT  605.36 0.0 605.92 976.68 ;
         LAYER MET4 ;
         RECT  29.44 0.0 30.0 976.68 ;
         LAYER MET4 ;
         RECT  750.72 0.0 751.28 976.68 ;
         LAYER MET3 ;
         RECT  0.0 353.28 142.24 353.84 ;
         LAYER MET4 ;
         RECT  791.2 0.0 791.76 976.68 ;
         LAYER MET4 ;
         RECT  189.52 12.88 190.08 976.68 ;
         LAYER MET4 ;
         RECT  49.68 0.0 50.24 976.68 ;
         LAYER MET4 ;
         RECT  290.72 0.0 291.28 976.68 ;
         LAYER MET4 ;
         RECT  892.4 0.0 892.96 976.68 ;
         LAYER MET3 ;
         RECT  0.0 169.28 117.4 169.84 ;
         LAYER MET3 ;
         RECT  0.0 671.6 899.4 672.16 ;
         LAYER MET3 ;
         RECT  0.0 44.16 899.4 44.72 ;
         LAYER MET3 ;
         RECT  755.32 329.36 899.4 329.92 ;
         LAYER MET3 ;
         RECT  0.0 655.04 899.4 655.6 ;
         LAYER MET3 ;
         RECT  0.0 531.76 899.4 532.32 ;
         LAYER MET4 ;
         RECT  631.12 0.0 631.68 976.68 ;
         LAYER MET3 ;
         RECT  733.24 86.48 899.4 87.04 ;
         LAYER MET3 ;
         RECT  0.0 136.16 117.4 136.72 ;
         LAYER MET3 ;
         RECT  731.4 820.64 899.4 821.2 ;
         LAYER MET3 ;
         RECT  0.0 940.24 899.4 940.8 ;
         LAYER MET4 ;
         RECT  176.64 0.0 177.2 976.68 ;
         LAYER MET3 ;
         RECT  0.0 493.12 899.4 493.68 ;
         LAYER MET4 ;
         RECT  369.84 0.0 370.4 976.68 ;
         LAYER MET4 ;
         RECT  467.36 0.0 467.92 976.68 ;
         LAYER MET3 ;
         RECT  733.24 907.12 899.4 907.68 ;
         LAYER MET4 ;
         RECT  728.64 0.0 729.2 976.68 ;
         LAYER MET3 ;
         RECT  0.0 266.8 117.4 267.36 ;
         LAYER MET3 ;
         RECT  0.0 461.84 899.4 462.4 ;
         LAYER MET3 ;
         RECT  0.0 437.92 899.4 438.48 ;
         LAYER MET3 ;
         RECT  0.0 960.48 860.76 961.04 ;
         LAYER MET4 ;
         RECT  46.0 0.0 46.56 976.68 ;
         LAYER MET4 ;
         RECT  529.92 0.0 530.48 976.68 ;
         LAYER MET3 ;
         RECT  0.0 783.84 899.4 784.4 ;
         LAYER MET4 ;
         RECT  358.8 6.44 359.36 976.68 ;
         LAYER MET4 ;
         RECT  340.4 0.0 340.96 976.68 ;
         LAYER MET4 ;
         RECT  480.24 0.0 480.8 976.68 ;
         LAYER MET3 ;
         RECT  780.16 110.4 899.4 110.96 ;
         LAYER MET4 ;
         RECT  638.48 0.0 639.04 976.68 ;
         LAYER MET3 ;
         RECT  731.4 559.36 899.4 559.92 ;
         LAYER MET3 ;
         RECT  0.0 927.36 740.24 927.92 ;
         LAYER MET3 ;
         RECT  733.24 160.08 899.4 160.64 ;
         LAYER MET4 ;
         RECT  450.8 0.0 451.36 11.6 ;
         LAYER MET3 ;
         RECT  716.68 439.76 899.4 440.32 ;
         LAYER MET4 ;
         RECT  156.4 12.88 156.96 976.68 ;
         LAYER MET3 ;
         RECT  0.0 794.88 160.64 795.44 ;
         LAYER MET3 ;
         RECT  0.0 964.16 821.2 964.72 ;
         LAYER MET4 ;
         RECT  472.88 0.0 473.44 976.68 ;
         LAYER MET4 ;
         RECT  296.24 0.0 296.8 976.68 ;
         LAYER MET3 ;
         RECT  0.0 861.12 899.4 861.68 ;
         LAYER MET3 ;
         RECT  417.68 14.72 899.4 15.28 ;
         LAYER MET4 ;
         RECT  281.52 0.0 282.08 11.6 ;
         LAYER MET4 ;
         RECT  138.0 0.0 138.56 976.68 ;
         LAYER MET4 ;
         RECT  890.56 0.0 891.12 976.68 ;
         LAYER MET3 ;
         RECT  0.0 152.72 899.4 153.28 ;
         LAYER MET3 ;
         RECT  716.68 489.44 899.4 490.0 ;
         LAYER MET3 ;
         RECT  0.0 607.2 899.4 607.76 ;
         LAYER MET4 ;
         RECT  682.64 0.0 683.2 976.68 ;
         LAYER MET3 ;
         RECT  0.0 410.32 899.4 410.88 ;
         LAYER MET3 ;
         RECT  0.0 572.24 899.4 572.8 ;
         LAYER MET3 ;
         RECT  0.0 171.12 117.4 171.68 ;
         LAYER MET3 ;
         RECT  0.0 730.48 899.4 731.04 ;
         LAYER MET3 ;
         RECT  755.32 776.48 899.4 777.04 ;
         LAYER MET3 ;
         RECT  0.0 206.08 117.4 206.64 ;
         LAYER MET4 ;
         RECT  414.0 0.0 414.56 976.68 ;
         LAYER MET3 ;
         RECT  0.0 954.96 179.04 955.52 ;
         LAYER MET3 ;
         RECT  716.68 165.6 899.4 166.16 ;
         LAYER MET3 ;
         RECT  0.0 252.08 899.4 252.64 ;
         LAYER MET3 ;
         RECT  716.68 364.32 899.4 364.88 ;
         LAYER MET3 ;
         RECT  0.0 816.96 899.4 817.52 ;
         LAYER MET4 ;
         RECT  412.16 0.0 412.72 976.68 ;
         LAYER MET4 ;
         RECT  632.96 0.0 633.52 976.68 ;
         LAYER MET3 ;
         RECT  0.0 932.88 899.4 933.44 ;
         LAYER MET4 ;
         RECT  546.48 0.0 547.04 976.68 ;
         LAYER MET3 ;
         RECT  0.0 770.96 162.48 771.52 ;
         LAYER MET3 ;
         RECT  817.88 84.64 899.4 85.2 ;
         LAYER MET3 ;
         RECT  716.68 342.24 899.4 342.8 ;
         LAYER MET3 ;
         RECT  0.0 460.0 899.4 460.56 ;
         LAYER MET4 ;
         RECT  408.48 0.0 409.04 976.68 ;
         LAYER MET4 ;
         RECT  16.56 0.0 17.12 976.68 ;
         LAYER MET3 ;
         RECT  733.24 447.12 899.4 447.68 ;
         LAYER MET3 ;
         RECT  0.0 507.84 899.4 508.4 ;
         LAYER MET4 ;
         RECT  171.12 0.0 171.68 976.68 ;
         LAYER MET4 ;
         RECT  406.64 0.0 407.2 976.68 ;
         LAYER MET4 ;
         RECT  496.8 0.0 497.36 976.68 ;
         LAYER MET4 ;
         RECT  747.04 0.0 747.6 976.68 ;
         LAYER MET3 ;
         RECT  0.0 478.4 142.24 478.96 ;
         LAYER MET4 ;
         RECT  141.68 0.0 142.24 976.68 ;
         LAYER MET3 ;
         RECT  0.0 149.04 160.64 149.6 ;
         LAYER MET3 ;
         RECT  0.0 690.0 177.2 690.56 ;
         LAYER MET3 ;
         RECT  733.24 708.4 899.4 708.96 ;
         LAYER MET4 ;
         RECT  23.92 0.0 24.48 976.68 ;
         LAYER MET4 ;
         RECT  257.6 0.0 258.16 976.68 ;
         LAYER MET3 ;
         RECT  0.0 58.88 7.0 59.44 ;
         LAYER MET4 ;
         RECT  237.36 0.0 237.92 976.68 ;
         LAYER MET3 ;
         RECT  733.24 322.0 899.4 322.56 ;
         LAYER MET4 ;
         RECT  55.2 0.0 55.76 976.68 ;
         LAYER MET3 ;
         RECT  0.0 307.28 899.4 307.84 ;
         LAYER MET3 ;
         RECT  0.0 647.68 899.4 648.24 ;
         LAYER MET3 ;
         RECT  0.0 754.4 899.4 754.96 ;
         LAYER MET4 ;
         RECT  382.72 0.0 383.28 9.76 ;
         LAYER MET3 ;
         RECT  0.0 638.48 177.2 639.04 ;
         LAYER MET4 ;
         RECT  684.48 0.0 685.04 976.68 ;
         LAYER MET4 ;
         RECT  555.68 0.0 556.24 976.68 ;
         LAYER MET4 ;
         RECT  38.64 0.0 39.2 976.68 ;
         LAYER MET3 ;
         RECT  733.24 745.2 899.4 745.76 ;
         LAYER MET3 ;
         RECT  0.0 609.04 162.48 609.6 ;
         LAYER MET4 ;
         RECT  526.24 0.0 526.8 976.68 ;
         LAYER MET3 ;
         RECT  755.32 627.44 899.4 628.0 ;
         LAYER MET4 ;
         RECT  250.24 0.0 250.8 976.68 ;
         LAYER MET3 ;
         RECT  0.0 583.28 160.64 583.84 ;
         LAYER MET4 ;
         RECT  798.56 0.0 799.12 976.68 ;
         LAYER MET3 ;
         RECT  780.16 246.56 899.4 247.12 ;
         LAYER MET3 ;
         RECT  93.84 294.4 899.4 294.96 ;
         LAYER MET3 ;
         RECT  716.68 465.52 899.4 466.08 ;
         LAYER MET4 ;
         RECT  443.44 0.0 444.0 976.68 ;
         LAYER MET4 ;
         RECT  448.96 0.0 449.52 962.88 ;
         LAYER MET3 ;
         RECT  895.16 958.64 899.4 959.2 ;
         LAYER MET3 ;
         RECT  0.0 150.88 899.4 151.44 ;
         LAYER MET3 ;
         RECT  0.0 688.16 177.2 688.72 ;
         LAYER MET3 ;
         RECT  0.0 831.68 160.64 832.24 ;
         LAYER MET4 ;
         RECT  191.36 0.0 191.92 976.68 ;
         LAYER MET4 ;
         RECT  307.28 0.0 307.84 976.68 ;
         LAYER MET4 ;
         RECT  851.92 0.0 852.48 976.68 ;
         LAYER MET3 ;
         RECT  0.0 160.08 160.64 160.64 ;
         LAYER MET4 ;
         RECT  723.12 0.0 723.68 976.68 ;
         LAYER MET3 ;
         RECT  0.0 121.44 117.4 122.0 ;
         LAYER MET3 ;
         RECT  0.0 526.24 899.4 526.8 ;
         LAYER MET3 ;
         RECT  0.0 782.0 160.64 782.56 ;
         LAYER MET3 ;
         RECT  0.0 721.28 899.4 721.84 ;
         LAYER MET3 ;
         RECT  0.0 717.6 899.4 718.16 ;
         LAYER MET4 ;
         RECT  172.96 12.88 173.52 976.68 ;
         LAYER MET4 ;
         RECT  312.8 0.0 313.36 962.88 ;
         LAYER MET4 ;
         RECT  390.08 0.0 390.64 976.68 ;
         LAYER MET3 ;
         RECT  716.68 739.68 899.4 740.24 ;
         LAYER MET3 ;
         RECT  45.08 27.6 899.4 28.16 ;
         LAYER MET3 ;
         RECT  0.0 653.2 899.4 653.76 ;
         LAYER MET4 ;
         RECT  60.72 0.0 61.28 976.68 ;
         LAYER MET4 ;
         RECT  621.92 0.0 622.48 976.68 ;
         LAYER MET4 ;
         RECT  693.68 0.0 694.24 976.68 ;
         LAYER MET4 ;
         RECT  228.16 0.0 228.72 976.68 ;
         LAYER MET4 ;
         RECT  557.52 0.0 558.08 976.68 ;
         LAYER MET3 ;
         RECT  0.0 693.68 899.4 694.24 ;
         LAYER MET3 ;
         RECT  0.0 822.48 899.4 823.04 ;
         LAYER MET3 ;
         RECT  0.0 217.12 177.2 217.68 ;
         LAYER MET3 ;
         RECT  780.16 209.76 899.4 210.32 ;
         LAYER MET4 ;
         RECT  1.84 0.0 2.4 54.84 ;
         LAYER MET4 ;
         RECT  785.68 0.0 786.24 976.68 ;
         LAYER MET3 ;
         RECT  0.0 894.24 160.64 894.8 ;
         LAYER MET4 ;
         RECT  651.36 0.0 651.92 962.88 ;
         LAYER MET3 ;
         RECT  716.68 215.28 899.4 215.84 ;
         LAYER MET3 ;
         RECT  0.0 776.48 142.24 777.04 ;
         LAYER MET3 ;
         RECT  0.0 741.52 899.4 742.08 ;
         LAYER MET3 ;
         RECT  0.0 594.32 899.4 594.88 ;
         LAYER MET4 ;
         RECT  40.48 0.0 41.04 976.68 ;
      END
   END gnd
   OBS
   LAYER  MET1 ;
      RECT  0.0 0.0 899.4 976.68 ;
   LAYER  MET2 ;
      RECT  0.0 0.0 899.4 976.68 ;
   LAYER  MET3 ;
      RECT  161.36 191.72 779.44 193.4 ;
      RECT  161.36 193.4 779.44 195.4 ;
      RECT  118.12 279.88 161.36 281.88 ;
      RECT  161.36 182.36 779.44 184.36 ;
      RECT  177.92 165.96 715.96 173.16 ;
      RECT  2.2 86.84 177.92 87.6 ;
      RECT  161.36 178.84 177.92 182.36 ;
      RECT  177.92 178.84 715.96 182.36 ;
      RECT  715.96 178.84 779.44 182.36 ;
      RECT  177.0 961.76 752.92 962.52 ;
      RECT  161.36 191.56 732.52 191.72 ;
      RECT  118.12 92.36 161.36 97.72 ;
      RECT  161.36 184.36 779.44 186.04 ;
      RECT  118.12 178.84 161.36 186.04 ;
      RECT  110.76 4.04 121.8 5.88 ;
      RECT  161.36 195.4 732.52 198.92 ;
      RECT  78.56 320.36 79.32 320.52 ;
      RECT  2.2 0.0 397.64 0.2 ;
      RECT  397.64 0.0 405.0 0.2 ;
      RECT  405.0 0.0 820.84 0.2 ;
      RECT  820.84 0.0 897.2 0.2 ;
      RECT  897.2 0.0 899.4 0.2 ;
      RECT  121.8 38.84 131.76 39.0 ;
      RECT  73.96 294.6 92.2 294.76 ;
      RECT  23.36 11.4 30.72 13.08 ;
      RECT  2.2 303.8 79.32 303.96 ;
      RECT  90.36 9.56 121.8 11.4 ;
      RECT  0.0 0.0 2.2 0.2 ;
      RECT  161.36 129.16 715.96 136.36 ;
      RECT  715.96 129.16 779.44 136.36 ;
      RECT  118.12 129.16 161.36 136.36 ;
      RECT  740.96 925.88 752.92 927.56 ;
      RECT  740.96 925.72 752.92 925.88 ;
      RECT  78.56 329.56 79.32 329.72 ;
      RECT  30.72 16.92 121.8 18.6 ;
      RECT  121.8 16.92 179.76 18.6 ;
      RECT  179.76 16.92 186.2 18.6 ;
      RECT  271.76 14.92 405.0 16.92 ;
      RECT  177.92 116.28 715.96 123.48 ;
      RECT  715.96 92.36 732.52 99.56 ;
      RECT  865.16 958.84 876.96 959.0 ;
      RECT  118.12 254.28 161.36 261.48 ;
      RECT  161.36 254.28 732.52 261.48 ;
      RECT  732.52 254.28 779.44 261.48 ;
      RECT  110.76 3.88 393.96 4.04 ;
      RECT  186.2 4.04 393.96 5.88 ;
      RECT  177.92 856.88 715.96 857.64 ;
      RECT  177.92 869.76 715.96 870.52 ;
      RECT  177.92 589.16 715.96 590.08 ;
      RECT  177.92 590.08 715.96 590.84 ;
      RECT  177.92 894.44 715.96 895.36 ;
      RECT  177.92 757.52 715.96 758.28 ;
      RECT  177.92 414.36 715.96 415.28 ;
      RECT  177.92 415.28 715.96 416.04 ;
      RECT  90.52 62.92 171.48 63.68 ;
      RECT  171.48 62.92 732.52 63.68 ;
      RECT  2.2 62.92 7.72 63.68 ;
      RECT  7.72 62.92 90.52 63.68 ;
      RECT  0.0 62.92 2.2 63.68 ;
      RECT  405.0 10.48 654.32 11.4 ;
      RECT  271.76 9.56 397.64 10.48 ;
      RECT  271.76 10.48 397.64 14.92 ;
      RECT  397.64 10.48 405.0 14.92 ;
      RECT  0.0 79.48 2.2 80.24 ;
      RECT  816.4 79.48 819.16 80.24 ;
      RECT  819.16 79.48 820.84 80.24 ;
      RECT  2.2 79.48 16.76 80.24 ;
      RECT  16.76 79.48 177.92 80.24 ;
      RECT  177.92 79.48 816.4 80.24 ;
      RECT  177.92 322.36 715.96 323.12 ;
      RECT  90.52 62.0 816.4 62.92 ;
      RECT  897.2 876.2 899.4 876.96 ;
      RECT  883.56 876.2 897.2 876.96 ;
      RECT  881.72 876.2 883.56 876.96 ;
      RECT  177.92 490.56 715.96 491.48 ;
      RECT  177.92 887.24 715.96 888.16 ;
      RECT  5.88 11.4 23.36 12.16 ;
      RECT  2.2 53.72 18.6 54.64 ;
      RECT  2.2 54.64 18.6 55.56 ;
      RECT  18.6 54.64 820.84 55.56 ;
      RECT  850.44 954.4 856.88 955.16 ;
      RECT  856.88 954.4 865.16 955.16 ;
      RECT  865.16 954.4 869.6 955.16 ;
      RECT  101.56 92.36 118.12 93.12 ;
      RECT  741.88 972.8 752.92 973.56 ;
      RECT  142.96 315.92 177.92 316.68 ;
      RECT  861.48 959.92 897.2 960.84 ;
      RECT  861.48 959.0 865.16 959.76 ;
      RECT  177.92 496.24 715.96 497.0 ;
      RECT  732.52 195.4 779.44 198.0 ;
      RECT  177.92 521.08 715.96 521.84 ;
      RECT  881.72 918.52 883.56 919.28 ;
      RECT  883.56 918.52 891.68 919.28 ;
      RECT  891.68 918.52 897.2 919.28 ;
      RECT  897.2 918.52 899.4 919.28 ;
      RECT  752.92 970.96 771.16 971.88 ;
      RECT  752.92 961.76 867.76 963.44 ;
      RECT  177.92 787.88 715.96 788.64 ;
      RECT  177.92 788.64 715.96 789.56 ;
      RECT  177.92 789.56 715.96 789.72 ;
      RECT  897.2 901.96 899.4 902.72 ;
      RECT  883.56 901.96 897.2 902.72 ;
      RECT  881.72 901.96 883.56 902.72 ;
      RECT  161.36 166.88 177.92 173.16 ;
      RECT  118.12 166.88 161.36 173.16 ;
      RECT  732.52 241.4 779.44 247.68 ;
      RECT  177.92 863.16 732.52 863.32 ;
      RECT  73.96 293.84 81.32 294.6 ;
      RECT  81.32 293.84 92.2 294.6 ;
      RECT  177.92 291.08 715.96 291.84 ;
      RECT  177.92 291.84 715.96 292.0 ;
      RECT  177.92 292.0 715.96 292.76 ;
      RECT  177.92 384.0 715.96 384.76 ;
      RECT  177.92 633.32 715.96 634.08 ;
      RECT  177.92 539.48 715.96 540.24 ;
      RECT  177.92 540.24 715.96 541.16 ;
      RECT  177.92 141.12 715.96 142.8 ;
      RECT  177.92 142.8 715.96 143.72 ;
      RECT  78.56 328.8 79.32 329.56 ;
      RECT  79.32 328.8 96.8 329.56 ;
      RECT  177.92 396.88 715.96 397.64 ;
      RECT  805.36 88.52 825.44 89.44 ;
      RECT  825.44 88.52 897.2 89.44 ;
      RECT  177.92 688.52 715.96 691.12 ;
      RECT  177.92 173.16 715.96 174.08 ;
      RECT  161.36 190.8 732.52 191.56 ;
      RECT  0.0 103.4 2.2 104.16 ;
      RECT  78.56 336.16 79.32 337.08 ;
      RECT  715.96 117.2 779.44 123.48 ;
      RECT  177.92 85.92 715.96 86.84 ;
      RECT  2.2 310.4 79.32 311.32 ;
      RECT  161.36 309.48 715.96 310.24 ;
      RECT  177.92 813.64 715.96 814.4 ;
      RECT  177.92 814.4 715.96 815.32 ;
      RECT  177.92 707.84 715.96 708.6 ;
      RECT  177.92 160.44 715.96 161.2 ;
      RECT  161.36 240.48 715.96 248.6 ;
      RECT  715.96 240.48 732.52 248.6 ;
      RECT  177.92 341.68 715.96 342.44 ;
      RECT  90.52 55.56 816.4 56.32 ;
      RECT  2.2 55.56 88.68 56.32 ;
      RECT  88.68 55.56 90.52 56.32 ;
      RECT  0.0 53.72 2.2 56.32 ;
      RECT  816.4 55.56 817.16 56.32 ;
      RECT  817.16 55.56 820.84 56.32 ;
      RECT  32.56 9.4 90.36 9.56 ;
      RECT  5.88 10.48 32.56 11.4 ;
      RECT  32.56 9.56 90.36 10.48 ;
      RECT  32.56 10.48 90.36 11.4 ;
      RECT  177.92 488.88 715.96 490.56 ;
      RECT  118.12 279.12 161.36 279.88 ;
      RECT  7.72 112.6 18.6 113.36 ;
      RECT  2.2 112.6 7.72 113.36 ;
      RECT  0.0 112.6 2.2 113.36 ;
      RECT  177.92 638.84 715.96 639.6 ;
      RECT  177.92 639.6 715.96 640.52 ;
      RECT  177.92 440.12 715.96 440.88 ;
      RECT  177.92 440.88 715.96 441.8 ;
      RECT  161.36 117.2 177.92 123.48 ;
      RECT  118.12 117.2 161.36 123.48 ;
      RECT  816.4 71.2 820.84 71.96 ;
      RECT  118.12 266.24 161.36 273.44 ;
      RECT  161.36 266.24 177.92 273.44 ;
      RECT  177.92 266.24 732.52 273.44 ;
      RECT  897.2 892.76 899.4 893.52 ;
      RECT  754.6 892.76 883.56 893.52 ;
      RECT  883.56 892.76 897.2 893.52 ;
      RECT  177.92 812.72 715.96 813.64 ;
      RECT  0.0 86.84 2.2 87.6 ;
      RECT  177.92 738.2 715.96 738.96 ;
      RECT  177.92 738.96 715.96 739.88 ;
      RECT  2.2 70.28 7.72 71.04 ;
      RECT  0.0 70.28 2.2 71.04 ;
      RECT  161.36 73.04 732.52 73.8 ;
      RECT  803.52 71.2 816.4 71.96 ;
      RECT  7.72 70.28 18.6 71.04 ;
      RECT  177.92 421.72 715.96 422.48 ;
      RECT  732.52 62.92 738.96 63.68 ;
      RECT  738.96 62.92 816.4 63.68 ;
      RECT  171.48 63.68 714.12 64.6 ;
      RECT  816.4 62.0 820.84 63.68 ;
      RECT  110.76 3.12 397.64 3.88 ;
      RECT  397.64 3.12 405.0 3.88 ;
      RECT  90.52 3.12 110.76 3.88 ;
      RECT  114.44 0.2 397.64 1.12 ;
      RECT  78.56 337.08 79.32 337.84 ;
      RECT  79.32 337.08 97.72 337.84 ;
      RECT  2.2 336.16 78.56 337.84 ;
      RECT  177.92 339.84 715.96 341.68 ;
      RECT  177.92 372.04 715.96 372.8 ;
      RECT  856.88 950.72 865.92 951.48 ;
      RECT  754.6 926.64 808.88 927.56 ;
      RECT  177.92 837.56 715.96 838.32 ;
      RECT  177.92 838.32 715.96 839.24 ;
      RECT  121.8 38.08 131.76 38.84 ;
      RECT  131.76 38.08 157.52 38.84 ;
      RECT  90.52 38.08 121.8 38.84 ;
      RECT  2.2 303.04 79.32 303.8 ;
      RECT  883.56 909.32 897.2 910.08 ;
      RECT  897.2 909.32 899.4 910.08 ;
      RECT  881.72 909.32 883.56 910.08 ;
      RECT  30.72 11.4 121.8 14.0 ;
      RECT  23.36 13.08 30.72 14.0 ;
      RECT  121.8 9.56 179.76 14.0 ;
      RECT  179.76 9.56 186.2 14.0 ;
      RECT  186.2 9.56 271.76 14.0 ;
      RECT  177.92 416.04 715.96 416.2 ;
      RECT  78.56 319.6 79.32 320.36 ;
      RECT  177.92 234.96 715.96 235.72 ;
      RECT  865.16 958.08 876.96 958.84 ;
      RECT  2.2 303.96 79.32 304.72 ;
      RECT  79.32 303.96 94.04 304.72 ;
      RECT  121.8 4.04 179.76 6.64 ;
      RECT  179.76 4.04 186.2 6.64 ;
      RECT  110.76 5.88 121.8 6.64 ;
      RECT  186.2 5.88 393.96 6.64 ;
      RECT  393.96 5.88 405.0 6.64 ;
      RECT  32.56 8.64 90.36 9.4 ;
      RECT  177.92 334.32 715.96 335.08 ;
      RECT  177.92 732.68 715.96 733.44 ;
      RECT  177.92 364.68 715.96 365.6 ;
      RECT  177.92 365.6 715.96 366.36 ;
      RECT  177.92 832.04 715.96 832.8 ;
      RECT  121.8 39.0 131.76 39.76 ;
      RECT  177.92 123.48 715.96 124.4 ;
      RECT  177.92 366.52 715.96 367.28 ;
      RECT  177.92 770.4 715.96 771.16 ;
      RECT  78.56 329.72 79.32 330.48 ;
      RECT  177.92 545.92 715.96 546.68 ;
      RECT  177.92 347.2 715.96 347.96 ;
      RECT  28.88 50.96 37.92 51.72 ;
      RECT  177.92 713.36 715.96 715.04 ;
      RECT  177.92 763.8 715.96 763.96 ;
      RECT  177.92 763.04 715.96 763.8 ;
      RECT  177.92 763.96 715.96 764.72 ;
      RECT  33.48 20.6 42.52 21.36 ;
      RECT  177.92 315.0 715.96 315.92 ;
      RECT  873.28 960.84 897.2 961.6 ;
      RECT  867.76 961.76 873.28 963.44 ;
      RECT  78.56 320.52 95.88 321.28 ;
      RECT  88.68 66.6 90.36 67.36 ;
      RECT  2.2 103.4 18.6 104.16 ;
      RECT  101.56 104.32 118.12 105.08 ;
      RECT  177.92 807.2 715.96 807.96 ;
      RECT  177.92 789.72 715.96 790.48 ;
      RECT  715.96 893.68 732.52 894.44 ;
      RECT  753.84 892.76 754.6 893.52 ;
      RECT  177.92 148.48 715.96 149.24 ;
      RECT  161.36 91.44 715.96 99.56 ;
      RECT  715.96 91.44 732.52 92.36 ;
      RECT  807.2 89.44 825.44 89.6 ;
      RECT  807.2 89.6 825.44 90.36 ;
      RECT  177.92 863.32 715.96 864.08 ;
      RECT  177.92 864.08 715.96 864.24 ;
      RECT  715.96 863.32 754.6 864.08 ;
      RECT  177.92 864.24 715.96 865.0 ;
      RECT  177.92 514.64 715.96 516.32 ;
      RECT  177.92 839.24 715.96 840.16 ;
      RECT  752.92 917.6 754.6 918.36 ;
      RECT  754.6 917.6 808.88 918.36 ;
      RECT  118.12 281.88 161.36 286.32 ;
      RECT  161.36 279.12 732.52 286.32 ;
      RECT  732.52 279.12 779.44 286.32 ;
      RECT  897.2 867.92 899.4 868.68 ;
      RECT  883.56 867.92 897.2 868.68 ;
      RECT  881.72 867.92 883.56 868.68 ;
      RECT  177.92 471.4 715.96 472.16 ;
      RECT  2.2 976.48 752.92 976.68 ;
      RECT  752.92 976.48 897.2 976.68 ;
      RECT  0.0 976.48 2.2 976.68 ;
      RECT  897.2 976.48 899.4 976.68 ;
      RECT  177.92 359.16 715.96 359.92 ;
      RECT  179.76 18.6 186.2 19.52 ;
      RECT  654.32 18.6 688.36 19.52 ;
      RECT  186.2 16.92 271.76 19.52 ;
      RECT  271.76 16.92 405.0 19.52 ;
      RECT  405.0 16.92 552.2 19.52 ;
      RECT  177.92 683.0 715.96 683.76 ;
      RECT  752.92 924.96 754.6 927.56 ;
      RECT  720.72 924.96 740.96 925.72 ;
      RECT  740.96 924.96 752.92 925.72 ;
      RECT  883.56 924.96 891.68 926.64 ;
      RECT  891.68 924.96 897.2 926.64 ;
      RECT  897.2 924.96 899.4 926.64 ;
      RECT  754.6 924.96 808.88 926.64 ;
      RECT  808.88 924.96 881.72 926.64 ;
      RECT  881.72 924.96 883.56 926.64 ;
      RECT  177.92 215.64 715.96 216.4 ;
      RECT  177.92 216.4 715.96 216.56 ;
      RECT  177.92 216.56 715.96 218.24 ;
      RECT  177.92 223.0 715.96 223.76 ;
      RECT  161.36 316.68 715.96 316.84 ;
      RECT  177.92 315.92 715.96 316.68 ;
      RECT  161.36 316.84 715.96 317.6 ;
      RECT  177.92 620.44 715.96 621.2 ;
      RECT  177.92 558.8 715.96 559.56 ;
      RECT  118.12 97.72 161.36 98.64 ;
      RECT  118.12 191.72 161.36 198.0 ;
      RECT  897.2 884.48 899.4 885.24 ;
      RECT  883.56 884.48 897.2 885.24 ;
      RECT  881.72 884.48 883.56 885.24 ;
      RECT  177.92 881.72 715.96 882.48 ;
      RECT  732.52 92.36 779.44 98.64 ;
      RECT  177.92 366.36 715.96 366.52 ;
      RECT  405.0 11.4 451.0 12.16 ;
      RECT  405.0 12.16 451.0 13.08 ;
      RECT  451.0 11.4 586.24 12.16 ;
      RECT  586.24 11.4 654.32 12.16 ;
      RECT  800.76 46.2 820.84 47.12 ;
      RECT  186.2 49.12 405.0 49.88 ;
      RECT  405.0 49.12 720.56 49.88 ;
      RECT  2.2 311.32 79.32 312.08 ;
      RECT  89.6 312.24 94.96 313.0 ;
      RECT  177.92 446.56 715.96 447.32 ;
      RECT  177.92 290.16 715.96 291.08 ;
      RECT  654.32 17.84 688.36 18.6 ;
      RECT  552.2 17.84 586.24 19.52 ;
      RECT  586.24 17.84 654.32 19.52 ;
      RECT  118.12 203.68 161.36 210.88 ;
      RECT  161.36 203.68 732.52 210.88 ;
      RECT  732.52 203.68 779.44 210.88 ;
      RECT  177.92 389.52 715.96 392.12 ;
      RECT  177.92 844.92 715.96 845.68 ;
      RECT  732.52 266.24 779.44 273.44 ;
      RECT  177.92 265.32 715.96 266.24 ;
      RECT  177.92 416.2 715.96 416.96 ;
      RECT  855.04 943.36 868.68 944.12 ;
      RECT  177.92 820.08 715.96 820.84 ;
      RECT  118.12 241.4 161.36 247.68 ;
      RECT  752.92 971.88 771.16 972.8 ;
      RECT  752.92 972.8 771.16 973.56 ;
      RECT  771.16 972.8 807.96 973.56 ;
      RECT  2.2 96.04 101.56 96.8 ;
      RECT  101.56 96.04 118.12 96.8 ;
      RECT  0.0 96.04 2.2 96.8 ;
      RECT  177.92 464.96 715.96 466.64 ;
      RECT  177.92 888.16 715.96 888.92 ;
      RECT  177.92 888.92 715.96 889.08 ;
      RECT  177.92 889.08 715.96 889.84 ;
      RECT  819.16 78.56 820.84 79.48 ;
      RECT  177.92 538.56 715.96 539.48 ;
      RECT  177.92 658.16 715.96 658.92 ;
      RECT  161.36 104.32 715.96 111.52 ;
      RECT  715.96 104.32 779.44 111.52 ;
      RECT  118.12 104.32 161.36 111.52 ;
      RECT  73.96 294.76 93.12 295.52 ;
      RECT  177.92 297.52 715.96 298.28 ;
      RECT  177.92 670.12 715.96 670.88 ;
      RECT  186.2 45.44 405.0 46.2 ;
      RECT  121.8 45.44 157.52 46.2 ;
      RECT  157.52 45.44 186.2 46.2 ;
      RECT  0.0 45.44 2.2 46.2 ;
      RECT  2.2 45.44 31.64 46.2 ;
      RECT  31.64 45.44 121.8 46.2 ;
      RECT  405.0 45.44 720.56 46.2 ;
      RECT  720.56 45.44 800.76 46.2 ;
      RECT  800.76 45.44 820.84 46.2 ;
      RECT  805.36 87.76 897.2 88.52 ;
      RECT  177.92 86.84 732.52 87.6 ;
      RECT  142.96 87.6 732.52 87.76 ;
      RECT  142.96 87.76 732.52 88.52 ;
      RECT  732.52 87.76 805.36 88.52 ;
      RECT  161.36 907.48 732.52 908.24 ;
      RECT  177.92 439.2 715.96 440.12 ;
      RECT  861.48 960.84 873.28 961.6 ;
      RECT  861.48 961.6 873.28 961.76 ;
      RECT  177.92 782.36 715.96 783.12 ;
      RECT  177.0 962.52 752.92 963.44 ;
      RECT  821.92 963.44 867.76 964.36 ;
      RECT  715.96 862.4 732.52 863.16 ;
      RECT  881.72 859.64 897.2 860.4 ;
      RECT  897.2 859.64 899.4 860.4 ;
      RECT  177.92 862.4 715.96 863.16 ;
      RECT  405.0 14.92 416.96 15.08 ;
      RECT  405.0 15.08 416.96 16.0 ;
      RECT  405.0 16.0 416.96 16.92 ;
      RECT  416.96 16.0 552.2 16.92 ;
      RECT  405.0 13.08 416.96 14.0 ;
      RECT  405.0 14.0 416.96 14.16 ;
      RECT  416.96 13.08 451.0 14.0 ;
      RECT  405.0 14.16 416.96 14.92 ;
      RECT  177.92 608.48 715.96 609.24 ;
      RECT  177.92 408.84 715.96 409.6 ;
      RECT  177.92 570.76 715.96 571.52 ;
      RECT  715.96 166.88 779.44 173.16 ;
      RECT  766.72 934.16 808.88 934.92 ;
      RECT  740.04 934.16 766.72 934.92 ;
      RECT  177.92 458.52 715.96 459.28 ;
      RECT  177.92 509.12 715.96 509.88 ;
      RECT  865.16 959.0 894.44 959.76 ;
      RECT  861.48 959.76 894.44 959.92 ;
      RECT  177.92 719.8 715.96 720.56 ;
      RECT  31.64 27.96 44.36 28.72 ;
      RECT  161.36 893.68 715.96 894.44 ;
      RECT  177.92 739.88 715.96 740.8 ;
      RECT  177.92 595.6 715.96 596.36 ;
   LAYER  MET4 ;
      RECT  211.96 14.0 213.64 19.52 ;
      RECT  211.96 19.52 213.64 974.48 ;
      RECT  160.44 2.2 162.12 5.72 ;
      RECT  211.96 12.32 213.64 14.0 ;
      RECT  447.48 963.6 449.16 974.48 ;
      RECT  0.0 0.0 0.2 2.2 ;
      RECT  0.0 2.2 0.2 55.56 ;
      RECT  0.0 55.56 0.2 976.68 ;
      RECT  819.16 2.2 821.0 45.28 ;
      RECT  861.48 959.92 863.16 974.48 ;
      RECT  210.12 2.2 211.8 5.72 ;
      RECT  278.2 963.6 279.88 974.48 ;
      RECT  342.6 2.2 344.28 5.72 ;
      RECT  769.48 970.96 771.16 974.48 ;
      RECT  359.16 2.2 360.84 5.72 ;
      RECT  0.2 55.56 2.04 113.36 ;
      RECT  178.68 14.0 180.52 19.52 ;
      RECT  178.68 10.48 180.52 14.0 ;
      RECT  292.92 2.2 294.6 5.72 ;
      RECT  188.96 5.88 189.72 12.16 ;
      RECT  271.76 5.88 272.52 14.0 ;
      RECT  271.76 14.0 272.52 15.84 ;
      RECT  349.04 14.16 349.8 19.52 ;
      RECT  653.56 10.48 654.32 19.52 ;
      RECT  246.92 14.0 247.68 15.84 ;
      RECT  246.92 15.84 247.68 19.52 ;
      RECT  246.92 10.48 247.68 14.0 ;
      RECT  585.48 17.84 586.24 19.52 ;
      RECT  585.48 14.16 586.24 17.84 ;
      RECT  404.24 5.88 405.0 10.48 ;
      RECT  404.24 10.48 405.0 12.16 ;
      RECT  404.24 12.16 405.0 14.0 ;
      RECT  404.24 14.0 405.0 19.52 ;
      RECT  484.28 16.0 485.04 19.52 ;
      RECT  143.88 2.2 144.64 5.72 ;
      RECT  155.84 5.88 156.6 12.16 ;
      RECT  315.0 12.32 315.76 14.0 ;
      RECT  315.0 14.0 315.76 15.84 ;
      RECT  315.0 15.84 315.76 19.52 ;
      RECT  304.88 5.88 305.64 14.0 ;
      RECT  304.88 14.0 305.64 15.84 ;
      RECT  516.48 963.6 517.24 974.48 ;
      RECT  205.52 5.88 206.28 14.0 ;
      RECT  616.76 963.6 617.52 974.48 ;
      RECT  619.52 17.84 620.28 19.52 ;
      RECT  276.36 2.2 277.12 5.72 ;
      RECT  382.16 10.48 382.92 14.0 ;
      RECT  381.24 963.6 382.16 974.48 ;
      RECT  382.16 14.0 382.92 963.6 ;
      RECT  382.16 963.6 382.92 974.48 ;
      RECT  518.32 12.32 519.08 14.0 ;
      RECT  518.32 14.0 519.08 19.52 ;
      RECT  899.2 2.2 899.4 859.64 ;
      RECT  899.2 859.64 899.4 959.92 ;
      RECT  899.2 0.0 899.4 2.2 ;
      RECT  255.2 5.88 255.96 12.16 ;
      RECT  550.52 963.6 551.44 974.48 ;
      RECT  551.44 16.0 552.2 963.6 ;
      RECT  551.44 963.6 552.2 974.48 ;
      RECT  338.0 5.88 338.76 14.0 ;
      RECT  338.0 14.0 338.76 15.84 ;
      RECT  338.0 15.84 338.76 17.68 ;
      RECT  354.56 5.88 355.32 14.0 ;
      RECT  821.0 2.2 821.76 45.28 ;
      RECT  821.0 45.28 821.76 71.04 ;
      RECT  321.44 5.88 322.2 12.16 ;
      RECT  288.32 5.88 289.08 12.32 ;
      RECT  288.32 12.32 289.08 14.0 ;
      RECT  260.72 2.2 261.48 5.72 ;
      RECT  280.96 12.32 281.72 14.0 ;
      RECT  280.96 14.0 281.72 15.84 ;
      RECT  280.96 15.84 281.72 19.52 ;
      RECT  387.68 10.48 388.44 12.16 ;
      RECT  387.68 5.88 388.44 10.48 ;
      RECT  222.08 5.88 222.84 12.16 ;
      RECT  650.8 963.6 651.56 974.48 ;
      RECT  416.2 14.16 416.96 19.52 ;
      RECT  194.48 2.2 195.24 5.72 ;
      RECT  687.6 17.84 688.36 19.52 ;
      RECT  244.16 2.2 244.92 5.72 ;
      RECT  899.2 974.48 899.4 976.68 ;
      RECT  899.2 959.92 899.4 974.48 ;
      RECT  898.28 859.64 899.2 925.72 ;
      RECT  246.0 963.6 246.76 974.48 ;
      RECT  177.92 14.0 178.68 19.52 ;
      RECT  177.92 19.52 178.68 974.48 ;
      RECT  177.92 2.2 178.68 5.88 ;
      RECT  177.92 5.88 178.68 10.48 ;
      RECT  177.92 10.48 178.68 14.0 ;
      RECT  371.12 5.88 371.88 14.0 ;
      RECT  371.12 14.0 371.88 17.68 ;
      RECT  172.4 5.88 173.16 12.16 ;
      RECT  238.64 5.88 239.4 14.0 ;
      RECT  450.24 14.0 451.0 19.52 ;
      RECT  450.24 12.32 451.0 14.0 ;
      RECT  226.68 2.2 227.44 5.72 ;
   END
END    sram_0rw1r1w_16_256_lapis20
END    LIBRARY
