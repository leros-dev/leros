VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO sram_1rw0r0w_16_512_lapis20
   CLASS BLOCK ;
   SIZE 682.28 BY 578.32 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER MET4 ;
         RECT  166.52 0.0 167.08 1.48 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER MET4 ;
         RECT  184.0 0.0 184.56 1.48 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER MET4 ;
         RECT  200.56 0.0 201.12 1.48 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER MET4 ;
         RECT  216.2 0.0 216.76 1.48 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER MET4 ;
         RECT  232.76 0.0 233.32 1.48 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER MET4 ;
         RECT  250.24 0.0 250.8 1.48 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER MET4 ;
         RECT  266.8 0.0 267.36 1.48 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER MET4 ;
         RECT  282.44 0.0 283.0 1.48 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER MET4 ;
         RECT  299.0 0.0 299.56 1.48 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER MET4 ;
         RECT  316.48 0.0 317.04 1.48 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER MET4 ;
         RECT  333.04 0.0 333.6 1.48 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER MET4 ;
         RECT  348.68 0.0 349.24 1.48 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER MET4 ;
         RECT  365.24 0.0 365.8 1.48 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER MET4 ;
         RECT  382.72 0.0 383.28 1.48 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER MET4 ;
         RECT  399.28 0.0 399.84 1.48 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER MET4 ;
         RECT  414.92 0.0 415.48 1.48 ;
      END
   END din0[15]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER MET4 ;
         RECT  117.76 0.0 118.32 1.48 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER MET4 ;
         RECT  134.32 0.0 134.88 1.48 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER MET4 ;
         RECT  149.96 0.0 150.52 1.48 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER MET3 ;
         RECT  0.0 230.0 1.48 230.56 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER MET3 ;
         RECT  0.0 239.2 1.48 239.76 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER MET3 ;
         RECT  0.0 246.56 1.48 247.12 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER MET3 ;
         RECT  0.0 254.84 1.48 255.4 ;
      END
   END addr0[6]
   PIN addr0[7]
      DIRECTION INPUT ;
      PORT
         LAYER MET3 ;
         RECT  0.0 263.12 1.48 263.68 ;
      END
   END addr0[7]
   PIN addr0[8]
      DIRECTION INPUT ;
      PORT
         LAYER MET3 ;
         RECT  0.0 271.4 1.48 271.96 ;
      END
   END addr0[8]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER MET3 ;
         RECT  0.0 32.2 1.48 32.76 ;
      END
   END csb0
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER MET3 ;
         RECT  0.0 42.32 1.48 42.88 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER MET4 ;
         RECT  37.72 0.0 38.28 1.48 ;
      END
   END clk0
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER MET4 ;
         RECT  188.6 0.0 189.16 1.48 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER MET4 ;
         RECT  218.96 0.0 219.52 1.48 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER MET4 ;
         RECT  249.32 0.0 249.88 1.48 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER MET4 ;
         RECT  279.68 0.0 280.24 1.48 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER MET4 ;
         RECT  309.12 0.0 309.68 1.48 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER MET4 ;
         RECT  340.4 0.0 340.96 1.48 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER MET4 ;
         RECT  370.76 0.0 371.32 1.48 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER MET4 ;
         RECT  402.04 0.0 402.6 1.48 ;
      END
   END dout0[7]
   PIN dout0[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER MET4 ;
         RECT  431.48 0.0 432.04 1.48 ;
      END
   END dout0[8]
   PIN dout0[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER MET4 ;
         RECT  461.84 0.0 462.4 1.48 ;
      END
   END dout0[9]
   PIN dout0[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER MET4 ;
         RECT  493.12 0.0 493.68 1.48 ;
      END
   END dout0[10]
   PIN dout0[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER MET4 ;
         RECT  523.48 0.0 524.04 1.48 ;
      END
   END dout0[11]
   PIN dout0[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER MET4 ;
         RECT  553.84 0.0 554.4 1.48 ;
      END
   END dout0[12]
   PIN dout0[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER MET4 ;
         RECT  584.2 0.0 584.76 1.48 ;
      END
   END dout0[13]
   PIN dout0[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER MET4 ;
         RECT  614.56 0.0 615.12 1.48 ;
      END
   END dout0[14]
   PIN dout0[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER MET3 ;
         RECT  680.8 44.16 682.28 44.72 ;
      END
   END dout0[15]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER MET3 ;
         RECT  0.0 175.72 122.92 176.28 ;
         LAYER MET3 ;
         RECT  0.0 241.96 86.12 242.52 ;
         LAYER MET3 ;
         RECT  0.0 218.04 122.92 218.6 ;
         LAYER MET4 ;
         RECT  177.56 0.0 178.12 5.16 ;
         LAYER MET3 ;
         RECT  0.0 30.36 682.28 30.92 ;
         LAYER MET3 ;
         RECT  0.0 247.48 682.28 248.04 ;
         LAYER MET3 ;
         RECT  0.0 234.6 682.28 235.16 ;
         LAYER MET3 ;
         RECT  0.0 159.16 682.28 159.72 ;
         LAYER MET3 ;
         RECT  0.0 547.4 682.28 547.96 ;
         LAYER MET4 ;
         RECT  34.04 0.0 34.6 578.32 ;
         LAYER MET3 ;
         RECT  0.0 293.48 180.88 294.04 ;
         LAYER MET4 ;
         RECT  205.16 0.0 205.72 578.32 ;
         LAYER MET4 ;
         RECT  381.8 0.0 382.36 578.32 ;
         LAYER MET3 ;
         RECT  178.48 254.84 682.28 255.4 ;
         LAYER MET3 ;
         RECT  0.0 280.6 180.88 281.16 ;
         LAYER MET3 ;
         RECT  0.0 109.48 682.28 110.04 ;
         LAYER MET3 ;
         RECT  0.0 212.52 122.92 213.08 ;
         LAYER MET4 ;
         RECT  372.6 0.0 373.16 12.52 ;
         LAYER MET4 ;
         RECT  679.88 0.0 680.44 578.32 ;
         LAYER MET3 ;
         RECT  0.0 479.32 682.28 479.88 ;
         LAYER MET4 ;
         RECT  83.72 0.0 84.28 578.32 ;
         LAYER MET3 ;
         RECT  19.32 67.16 682.28 67.72 ;
         LAYER MET4 ;
         RECT  13.8 0.0 14.36 578.32 ;
         LAYER MET4 ;
         RECT  356.04 0.0 356.6 578.32 ;
         LAYER MET3 ;
         RECT  0.0 194.12 180.88 194.68 ;
         LAYER MET3 ;
         RECT  646.76 34.04 682.28 34.6 ;
         LAYER MET4 ;
         RECT  302.68 0.0 303.24 578.32 ;
         LAYER MET3 ;
         RECT  0.0 52.44 119.24 53.0 ;
         LAYER MET3 ;
         RECT  0.0 2.76 95.32 3.32 ;
         LAYER MET3 ;
         RECT  0.0 576.84 682.28 577.4 ;
         LAYER MET3 ;
         RECT  0.0 81.88 682.28 82.44 ;
         LAYER MET3 ;
         RECT  0.0 444.36 180.88 444.92 ;
         LAYER MET4 ;
         RECT  624.68 0.0 625.24 578.32 ;
         LAYER MET4 ;
         RECT  398.36 0.0 398.92 578.32 ;
         LAYER MET4 ;
         RECT  164.68 0.0 165.24 578.32 ;
         LAYER MET3 ;
         RECT  0.0 391.0 682.28 391.56 ;
         LAYER MET3 ;
         RECT  178.48 541.88 682.28 542.44 ;
         LAYER MET4 ;
         RECT  345.0 0.0 345.56 578.32 ;
         LAYER MET4 ;
         RECT  76.36 0.0 76.92 578.32 ;
         LAYER MET3 ;
         RECT  178.48 240.12 682.28 240.68 ;
         LAYER MET3 ;
         RECT  0.0 363.4 682.28 363.96 ;
         LAYER MET4 ;
         RECT  667.0 0.0 667.56 578.32 ;
         LAYER MET3 ;
         RECT  0.0 127.88 122.92 128.44 ;
         LAYER MET4 ;
         RECT  597.08 0.0 597.64 578.32 ;
         LAYER MET4 ;
         RECT  311.88 0.0 312.44 12.52 ;
         LAYER MET3 ;
         RECT  0.0 514.28 682.28 514.84 ;
         LAYER MET3 ;
         RECT  0.0 140.76 106.36 141.32 ;
         LAYER MET3 ;
         RECT  0.0 113.16 122.92 113.72 ;
         LAYER MET3 ;
         RECT  0.0 337.64 180.88 338.2 ;
         LAYER MET3 ;
         RECT  0.0 405.72 682.28 406.28 ;
         LAYER MET4 ;
         RECT  337.64 0.0 338.2 578.32 ;
         LAYER MET3 ;
         RECT  647.68 24.84 682.28 25.4 ;
         LAYER MET3 ;
         RECT  50.6 39.56 682.28 40.12 ;
         LAYER MET4 ;
         RECT  326.6 13.8 327.16 578.32 ;
         LAYER MET4 ;
         RECT  644.92 0.0 645.48 578.32 ;
         LAYER MET3 ;
         RECT  0.0 551.08 682.28 551.64 ;
         LAYER MET3 ;
         RECT  0.0 396.52 682.28 397.08 ;
         LAYER MET4 ;
         RECT  506.92 0.0 507.48 578.32 ;
         LAYER MET4 ;
         RECT  80.04 0.0 80.6 578.32 ;
         LAYER MET3 ;
         RECT  0.0 569.48 147.76 570.04 ;
         LAYER MET3 ;
         RECT  0.0 359.72 682.28 360.28 ;
         LAYER MET4 ;
         RECT  339.48 0.0 340.04 578.32 ;
         LAYER MET3 ;
         RECT  125.12 207.0 682.28 207.56 ;
         LAYER MET4 ;
         RECT  392.84 0.0 393.4 5.16 ;
         LAYER MET4 ;
         RECT  457.24 0.0 457.8 578.32 ;
         LAYER MET4 ;
         RECT  433.32 26.68 433.88 578.32 ;
         LAYER MET3 ;
         RECT  0.0 427.8 682.28 428.36 ;
         LAYER MET4 ;
         RECT  668.84 0.0 669.4 578.32 ;
         LAYER MET3 ;
         RECT  0.0 466.44 180.88 467.0 ;
         LAYER MET3 ;
         RECT  19.32 116.84 682.28 117.4 ;
         LAYER MET4 ;
         RECT  442.52 0.0 443.08 578.32 ;
         LAYER MET4 ;
         RECT  497.72 0.0 498.28 578.32 ;
         LAYER MET4 ;
         RECT  357.88 0.0 358.44 578.32 ;
         LAYER MET3 ;
         RECT  0.0 339.48 682.28 340.04 ;
         LAYER MET4 ;
         RECT  264.04 0.0 264.6 578.32 ;
         LAYER MET3 ;
         RECT  178.48 341.32 682.28 341.88 ;
         LAYER MET3 ;
         RECT  0.0 448.04 682.28 448.6 ;
         LAYER MET3 ;
         RECT  178.48 383.64 682.28 384.2 ;
         LAYER MET4 ;
         RECT  214.36 0.0 214.92 578.32 ;
         LAYER MET4 ;
         RECT  545.56 0.0 546.12 578.32 ;
         LAYER MET3 ;
         RECT  0.0 429.64 180.88 430.2 ;
         LAYER MET4 ;
         RECT  179.4 0.0 179.96 578.32 ;
         LAYER MET4 ;
         RECT  460.92 0.0 461.48 578.32 ;
         LAYER MET4 ;
         RECT  466.44 0.0 467.0 578.32 ;
         LAYER MET3 ;
         RECT  0.0 402.04 180.88 402.6 ;
         LAYER MET3 ;
         RECT  0.0 63.48 682.28 64.04 ;
         LAYER MET3 ;
         RECT  178.48 111.32 682.28 111.88 ;
         LAYER MET3 ;
         RECT  132.48 69.0 682.28 69.56 ;
         LAYER MET3 ;
         RECT  0.0 173.88 682.28 174.44 ;
         LAYER MET3 ;
         RECT  178.48 556.6 682.28 557.16 ;
         LAYER MET3 ;
         RECT  178.48 470.12 682.28 470.68 ;
         LAYER MET4 ;
         RECT  23.0 0.0 23.56 578.32 ;
         LAYER MET4 ;
         RECT  65.32 0.0 65.88 578.32 ;
         LAYER MET4 ;
         RECT  516.12 0.0 516.68 578.32 ;
         LAYER MET4 ;
         RECT  52.44 0.0 53.0 578.32 ;
         LAYER MET3 ;
         RECT  0.0 433.32 682.28 433.88 ;
         LAYER MET3 ;
         RECT  0.0 411.24 682.28 411.8 ;
         LAYER MET3 ;
         RECT  0.0 503.24 682.28 503.8 ;
         LAYER MET3 ;
         RECT  0.0 17.48 425.6 18.04 ;
         LAYER MET4 ;
         RECT  468.28 0.0 468.84 578.32 ;
         LAYER MET4 ;
         RECT  621.0 0.0 621.56 578.32 ;
         LAYER MET3 ;
         RECT  178.48 368.92 682.28 369.48 ;
         LAYER MET3 ;
         RECT  0.0 94.76 682.28 95.32 ;
         LAYER MET4 ;
         RECT  91.08 0.0 91.64 578.32 ;
         LAYER MET4 ;
         RECT  335.8 0.0 336.36 578.32 ;
         LAYER MET4 ;
         RECT  350.52 0.0 351.08 578.32 ;
         LAYER MET4 ;
         RECT  0.92 0.0 1.48 84.28 ;
         LAYER MET3 ;
         RECT  0.0 328.44 682.28 329.0 ;
         LAYER MET3 ;
         RECT  178.48 153.64 682.28 154.2 ;
         LAYER MET4 ;
         RECT  287.96 0.0 288.52 578.32 ;
         LAYER MET3 ;
         RECT  89.24 276.92 682.28 277.48 ;
         LAYER MET4 ;
         RECT  229.08 0.0 229.64 578.32 ;
         LAYER MET3 ;
         RECT  0.0 315.56 180.88 316.12 ;
         LAYER MET3 ;
         RECT  646.76 43.24 682.28 43.8 ;
         LAYER MET3 ;
         RECT  0.0 267.72 682.28 268.28 ;
         LAYER MET3 ;
         RECT  0.0 43.24 25.4 43.8 ;
         LAYER MET3 ;
         RECT  0.0 57.96 95.32 58.52 ;
         LAYER MET4 ;
         RECT  184.92 0.0 185.48 578.32 ;
         LAYER MET4 ;
         RECT  433.32 0.0 433.88 14.36 ;
         LAYER MET3 ;
         RECT  0.0 365.24 180.88 365.8 ;
         LAYER MET4 ;
         RECT  359.72 0.0 360.28 5.16 ;
         LAYER MET4 ;
         RECT  464.6 0.0 465.16 12.52 ;
         LAYER MET4 ;
         RECT  192.28 0.0 192.84 578.32 ;
         LAYER MET4 ;
         RECT  525.32 26.68 525.88 578.32 ;
         LAYER MET3 ;
         RECT  0.0 506.92 682.28 507.48 ;
         LAYER MET3 ;
         RECT  96.6 28.52 682.28 29.08 ;
         LAYER MET4 ;
         RECT  317.4 0.0 317.96 578.32 ;
         LAYER MET3 ;
         RECT  0.0 516.12 180.88 516.68 ;
         LAYER MET4 ;
         RECT  291.64 0.0 292.2 578.32 ;
         LAYER MET3 ;
         RECT  0.0 442.52 682.28 443.08 ;
         LAYER MET4 ;
         RECT  144.44 0.0 145.0 578.32 ;
         LAYER MET4 ;
         RECT  470.12 0.0 470.68 578.32 ;
         LAYER MET4 ;
         RECT  655.96 0.0 656.52 578.32 ;
         LAYER MET3 ;
         RECT  0.0 357.88 180.88 358.44 ;
         LAYER MET4 ;
         RECT  501.4 0.0 501.96 578.32 ;
         LAYER MET3 ;
         RECT  0.0 210.68 106.36 211.24 ;
         LAYER MET3 ;
         RECT  0.0 260.36 682.28 260.92 ;
         LAYER MET4 ;
         RECT  604.44 0.0 605.0 578.32 ;
         LAYER MET3 ;
         RECT  0.0 462.76 682.28 463.32 ;
         LAYER MET3 ;
         RECT  0.0 486.68 180.88 487.24 ;
         LAYER MET3 ;
         RECT  0.0 354.2 147.76 354.76 ;
         LAYER MET4 ;
         RECT  661.48 0.0 662.04 578.32 ;
         LAYER MET4 ;
         RECT  260.36 0.0 260.92 5.16 ;
         LAYER MET3 ;
         RECT  125.12 170.2 682.28 170.76 ;
         LAYER MET4 ;
         RECT  449.88 0.0 450.44 578.32 ;
         LAYER MET3 ;
         RECT  0.0 24.84 190.08 25.4 ;
         LAYER MET3 ;
         RECT  179.4 65.32 682.28 65.88 ;
         LAYER MET3 ;
         RECT  0.0 398.36 147.76 398.92 ;
         LAYER MET3 ;
         RECT  0.0 437.0 180.88 437.56 ;
         LAYER MET3 ;
         RECT  0.0 389.16 682.28 389.72 ;
         LAYER MET3 ;
         RECT  0.0 481.16 180.88 481.72 ;
         LAYER MET4 ;
         RECT  378.12 0.0 378.68 578.32 ;
         LAYER MET4 ;
         RECT  199.64 6.44 200.2 578.32 ;
         LAYER MET4 ;
         RECT  448.04 0.0 448.6 578.32 ;
         LAYER MET3 ;
         RECT  0.0 201.48 180.88 202.04 ;
         LAYER MET4 ;
         RECT  249.32 45.08 249.88 578.32 ;
         LAYER MET3 ;
         RECT  134.32 175.72 682.28 176.28 ;
         LAYER MET4 ;
         RECT  278.76 0.0 279.32 578.32 ;
         LAYER MET3 ;
         RECT  125.12 162.84 682.28 163.4 ;
         LAYER MET3 ;
         RECT  0.0 92.92 95.32 93.48 ;
         LAYER MET3 ;
         RECT  647.68 17.48 682.28 18.04 ;
         LAYER MET3 ;
         RECT  0.0 225.4 86.12 225.96 ;
         LAYER MET4 ;
         RECT  43.24 0.0 43.8 578.32 ;
         LAYER MET4 ;
         RECT  251.16 0.0 251.72 10.68 ;
         LAYER MET4 ;
         RECT  473.8 0.0 474.36 578.32 ;
         LAYER MET3 ;
         RECT  0.0 562.12 682.28 562.68 ;
         LAYER MET3 ;
         RECT  0.0 162.84 122.92 163.4 ;
         LAYER MET4 ;
         RECT  582.36 0.0 582.92 578.32 ;
         LAYER MET4 ;
         RECT  313.72 0.0 314.28 578.32 ;
         LAYER MET4 ;
         RECT  414.92 6.44 415.48 578.32 ;
         LAYER MET4 ;
         RECT  492.2 45.08 492.76 578.32 ;
         LAYER MET4 ;
         RECT  98.44 0.0 99.0 578.32 ;
         LAYER MET4 ;
         RECT  481.16 0.0 481.72 578.32 ;
         LAYER MET4 ;
         RECT  269.56 0.0 270.12 578.32 ;
         LAYER MET4 ;
         RECT  54.28 0.0 54.84 578.32 ;
         LAYER MET4 ;
         RECT  295.32 0.0 295.88 578.32 ;
         LAYER MET3 ;
         RECT  0.0 484.84 147.76 485.4 ;
         LAYER MET4 ;
         RECT  35.88 0.0 36.44 578.32 ;
         LAYER MET4 ;
         RECT  674.36 0.0 674.92 578.32 ;
         LAYER MET3 ;
         RECT  0.0 41.4 5.16 41.96 ;
         LAYER MET4 ;
         RECT  107.64 0.0 108.2 578.32 ;
         LAYER MET4 ;
         RECT  271.4 0.0 271.96 578.32 ;
         LAYER MET4 ;
         RECT  403.88 0.0 404.44 10.68 ;
         LAYER MET3 ;
         RECT  0.0 295.32 682.28 295.88 ;
         LAYER MET4 ;
         RECT  21.16 0.0 21.72 578.32 ;
         LAYER MET3 ;
         RECT  46.92 48.76 682.28 49.32 ;
         LAYER MET4 ;
         RECT  512.44 0.0 513.0 578.32 ;
         LAYER MET4 ;
         RECT  210.68 13.8 211.24 578.32 ;
         LAYER MET3 ;
         RECT  0.0 264.04 83.36 264.6 ;
         LAYER MET4 ;
         RECT  188.6 45.08 189.16 578.32 ;
         LAYER MET4 ;
         RECT  6.44 0.0 7.0 578.32 ;
         LAYER MET4 ;
         RECT  102.12 0.0 102.68 578.32 ;
         LAYER MET3 ;
         RECT  0.0 414.92 180.88 415.48 ;
         LAYER MET3 ;
         RECT  0.0 453.56 682.28 454.12 ;
         LAYER MET4 ;
         RECT  208.84 0.0 209.4 578.32 ;
         LAYER MET3 ;
         RECT  0.0 492.2 682.28 492.76 ;
         LAYER MET3 ;
         RECT  0.0 76.36 95.32 76.92 ;
         LAYER MET4 ;
         RECT  159.16 0.0 159.72 578.32 ;
         LAYER MET4 ;
         RECT  437.0 0.0 437.56 578.32 ;
         LAYER MET3 ;
         RECT  178.48 168.36 682.28 168.92 ;
         LAYER MET3 ;
         RECT  0.0 205.16 122.92 205.72 ;
         LAYER MET3 ;
         RECT  0.0 282.44 147.76 283.0 ;
         LAYER MET4 ;
         RECT  622.84 0.0 623.4 578.32 ;
         LAYER MET4 ;
         RECT  368.92 0.0 369.48 578.32 ;
         LAYER MET4 ;
         RECT  464.6 26.68 465.16 578.32 ;
         LAYER MET3 ;
         RECT  0.0 87.4 7.0 87.96 ;
         LAYER MET4 ;
         RECT  639.4 0.0 639.96 578.32 ;
         LAYER MET4 ;
         RECT  659.64 0.0 660.2 578.32 ;
         LAYER MET3 ;
         RECT  0.0 26.68 682.28 27.24 ;
         LAYER MET3 ;
         RECT  0.0 372.6 180.88 373.16 ;
         LAYER MET3 ;
         RECT  178.48 140.76 682.28 141.32 ;
         LAYER MET4 ;
         RECT  602.6 0.0 603.16 578.32 ;
         LAYER MET4 ;
         RECT  646.76 0.0 647.32 16.2 ;
         LAYER MET4 ;
         RECT  676.2 0.0 676.76 578.32 ;
         LAYER MET4 ;
         RECT  562.12 0.0 562.68 578.32 ;
         LAYER MET4 ;
         RECT  148.12 0.0 148.68 578.32 ;
         LAYER MET4 ;
         RECT  643.08 0.0 643.64 578.32 ;
         LAYER MET4 ;
         RECT  116.84 0.0 117.4 578.32 ;
         LAYER MET4 ;
         RECT  166.52 6.44 167.08 578.32 ;
         LAYER MET4 ;
         RECT  422.28 0.0 422.84 578.32 ;
         LAYER MET3 ;
         RECT  0.0 379.96 180.88 380.52 ;
         LAYER MET3 ;
         RECT  0.0 424.12 180.88 424.68 ;
         LAYER MET4 ;
         RECT  541.88 0.0 542.44 578.32 ;
         LAYER MET4 ;
         RECT  554.76 0.0 555.32 12.52 ;
         LAYER MET3 ;
         RECT  0.0 164.68 122.92 165.24 ;
         LAYER MET3 ;
         RECT  0.0 80.04 27.24 80.6 ;
         LAYER MET4 ;
         RECT  459.08 0.0 459.64 578.32 ;
         LAYER MET4 ;
         RECT  315.56 0.0 316.12 578.32 ;
         LAYER MET4 ;
         RECT  201.48 0.0 202.04 578.32 ;
         LAYER MET4 ;
         RECT  477.48 0.0 478.04 578.32 ;
         LAYER MET3 ;
         RECT  138.0 218.04 682.28 218.6 ;
         LAYER MET3 ;
         RECT  0.0 138.92 682.28 139.48 ;
         LAYER MET3 ;
         RECT  0.0 333.96 682.28 334.52 ;
         LAYER MET4 ;
         RECT  0.92 135.24 1.48 578.32 ;
         LAYER MET4 ;
         RECT  402.04 45.08 402.6 578.32 ;
         LAYER MET4 ;
         RECT  565.8 0.0 566.36 578.32 ;
         LAYER MET4 ;
         RECT  615.48 26.68 616.04 578.32 ;
         LAYER MET4 ;
         RECT  617.32 0.0 617.88 578.32 ;
         LAYER MET3 ;
         RECT  0.0 345.0 682.28 345.56 ;
         LAYER MET4 ;
         RECT  416.76 0.0 417.32 578.32 ;
         LAYER MET4 ;
         RECT  155.48 0.0 156.04 578.32 ;
         LAYER MET4 ;
         RECT  352.36 0.0 352.92 578.32 ;
         LAYER MET4 ;
         RECT  258.52 0.0 259.08 578.32 ;
         LAYER MET4 ;
         RECT  678.04 0.0 678.6 578.32 ;
         LAYER MET4 ;
         RECT  425.96 0.0 426.52 5.16 ;
         LAYER MET3 ;
         RECT  0.0 321.08 682.28 321.64 ;
         LAYER MET4 ;
         RECT  554.76 26.68 555.32 578.32 ;
         LAYER MET4 ;
         RECT  635.72 0.0 636.28 578.32 ;
         LAYER MET4 ;
         RECT  346.84 0.0 347.4 578.32 ;
         LAYER MET4 ;
         RECT  32.2 0.0 32.76 578.32 ;
         LAYER MET4 ;
         RECT  453.56 0.0 454.12 578.32 ;
         LAYER MET3 ;
         RECT  0.0 249.32 682.28 249.88 ;
         LAYER MET4 ;
         RECT  587.88 0.0 588.44 578.32 ;
         LAYER MET3 ;
         RECT  0.0 457.24 682.28 457.8 ;
         LAYER MET4 ;
         RECT  195.96 0.0 196.52 578.32 ;
         LAYER MET4 ;
         RECT  322.92 0.0 323.48 578.32 ;
         LAYER MET3 ;
         RECT  0.0 179.4 122.92 179.96 ;
         LAYER MET4 ;
         RECT  149.96 6.44 150.52 578.32 ;
         LAYER MET4 ;
         RECT  424.12 0.0 424.68 578.32 ;
         LAYER MET4 ;
         RECT  584.2 45.08 584.76 578.32 ;
         LAYER MET3 ;
         RECT  0.0 157.32 122.92 157.88 ;
         LAYER MET3 ;
         RECT  0.0 310.04 682.28 310.6 ;
         LAYER MET4 ;
         RECT  573.16 0.0 573.72 578.32 ;
         LAYER MET4 ;
         RECT  153.64 0.0 154.2 578.32 ;
         LAYER MET3 ;
         RECT  0.0 341.32 147.76 341.88 ;
         LAYER MET4 ;
         RECT  41.4 0.0 41.96 578.32 ;
         LAYER MET4 ;
         RECT  126.04 0.0 126.6 578.32 ;
         LAYER MET4 ;
         RECT  218.04 0.0 218.6 578.32 ;
         LAYER MET4 ;
         RECT  392.84 17.48 393.4 578.32 ;
         LAYER MET3 ;
         RECT  0.0 61.64 93.48 62.2 ;
         LAYER MET3 ;
         RECT  44.16 41.4 682.28 41.96 ;
         LAYER MET3 ;
         RECT  125.12 155.48 682.28 156.04 ;
         LAYER MET3 ;
         RECT  178.48 455.4 682.28 455.96 ;
         LAYER MET3 ;
         RECT  0.0 229.08 78.76 229.64 ;
         LAYER MET3 ;
         RECT  0.0 416.76 682.28 417.32 ;
         LAYER MET4 ;
         RECT  276.92 0.0 277.48 5.16 ;
         LAYER MET4 ;
         RECT  418.6 0.0 419.16 578.32 ;
         LAYER MET4 ;
         RECT  304.52 0.0 305.08 578.32 ;
         LAYER MET4 ;
         RECT  328.44 0.0 329.0 578.32 ;
         LAYER MET4 ;
         RECT  615.48 0.0 616.04 10.68 ;
         LAYER MET4 ;
         RECT  111.32 0.0 111.88 578.32 ;
         LAYER MET4 ;
         RECT  236.44 0.0 237.0 578.32 ;
         LAYER MET4 ;
         RECT  170.2 0.0 170.76 578.32 ;
         LAYER MET3 ;
         RECT  0.0 475.64 682.28 476.2 ;
         LAYER MET3 ;
         RECT  0.0 48.76 30.0 49.32 ;
         LAYER MET3 ;
         RECT  0.0 258.52 86.12 259.08 ;
         LAYER MET3 ;
         RECT  0.0 418.6 682.28 419.16 ;
         LAYER MET4 ;
         RECT  586.04 26.68 586.6 578.32 ;
         LAYER MET4 ;
         RECT  657.8 0.0 658.36 578.32 ;
         LAYER MET3 ;
         RECT  0.0 166.52 682.28 167.08 ;
         LAYER MET4 ;
         RECT  19.32 0.0 19.88 578.32 ;
         LAYER MET3 ;
         RECT  178.48 197.8 682.28 198.36 ;
         LAYER MET3 ;
         RECT  0.0 440.68 147.76 441.24 ;
         LAYER MET4 ;
         RECT  633.88 0.0 634.44 578.32 ;
         LAYER MET3 ;
         RECT  0.0 575.0 682.28 575.56 ;
         LAYER MET3 ;
         RECT  0.0 297.16 147.76 297.72 ;
         LAYER MET3 ;
         RECT  0.0 346.84 682.28 347.4 ;
         LAYER MET4 ;
         RECT  50.6 0.0 51.16 578.32 ;
         LAYER MET4 ;
         RECT  600.76 0.0 601.32 578.32 ;
         LAYER MET3 ;
         RECT  0.0 387.32 180.88 387.88 ;
         LAYER MET3 ;
         RECT  556.6 13.8 682.28 14.36 ;
         LAYER MET3 ;
         RECT  0.0 6.44 177.2 7.0 ;
         LAYER MET3 ;
         RECT  0.0 311.88 147.76 312.44 ;
         LAYER MET4 ;
         RECT  232.76 6.44 233.32 578.32 ;
         LAYER MET3 ;
         RECT  0.0 308.2 180.88 308.76 ;
         LAYER MET3 ;
         RECT  0.0 403.88 682.28 404.44 ;
         LAYER MET3 ;
         RECT  0.0 65.32 95.32 65.88 ;
         LAYER MET3 ;
         RECT  0.0 170.2 122.92 170.76 ;
         LAYER MET3 ;
         RECT  0.0 383.64 147.76 384.2 ;
         LAYER MET4 ;
         RECT  197.8 0.0 198.36 578.32 ;
         LAYER MET4 ;
         RECT  471.96 0.0 472.52 578.32 ;
         LAYER MET3 ;
         RECT  0.0 151.8 682.28 152.36 ;
         LAYER MET4 ;
         RECT  505.08 0.0 505.64 578.32 ;
         LAYER MET4 ;
         RECT  558.44 0.0 559.0 578.32 ;
         LAYER MET4 ;
         RECT  46.92 0.0 47.48 578.32 ;
         LAYER MET4 ;
         RECT  379.96 0.0 380.52 578.32 ;
         LAYER MET4 ;
         RECT  534.52 0.0 535.08 578.32 ;
         LAYER MET3 ;
         RECT  128.8 118.68 682.28 119.24 ;
         LAYER MET4 ;
         RECT  186.76 0.0 187.32 578.32 ;
         LAYER MET3 ;
         RECT  0.0 98.44 179.04 99.0 ;
         LAYER MET3 ;
         RECT  0.0 409.4 180.88 409.96 ;
         LAYER MET3 ;
         RECT  0.0 203.32 682.28 203.88 ;
         LAYER MET4 ;
         RECT  372.6 26.68 373.16 578.32 ;
         LAYER MET3 ;
         RECT  0.0 510.6 682.28 511.16 ;
         LAYER MET3 ;
         RECT  0.0 545.56 180.88 546.12 ;
         LAYER MET4 ;
         RECT  138.92 0.0 139.48 578.32 ;
         LAYER MET3 ;
         RECT  0.0 10.12 682.28 10.68 ;
         LAYER MET3 ;
         RECT  0.0 192.28 682.28 192.84 ;
         LAYER MET4 ;
         RECT  293.48 0.0 294.04 5.16 ;
         LAYER MET4 ;
         RECT  234.6 0.0 235.16 578.32 ;
         LAYER MET3 ;
         RECT  0.0 265.88 180.88 266.44 ;
         LAYER MET3 ;
         RECT  178.48 569.48 682.28 570.04 ;
         LAYER MET4 ;
         RECT  495.88 0.0 496.44 578.32 ;
         LAYER MET3 ;
         RECT  0.0 50.6 682.28 51.16 ;
         LAYER MET4 ;
         RECT  521.64 0.0 522.2 578.32 ;
         LAYER MET3 ;
         RECT  0.0 37.72 682.28 38.28 ;
         LAYER MET4 ;
         RECT  100.28 0.0 100.84 578.32 ;
         LAYER MET4 ;
         RECT  462.76 0.0 463.32 578.32 ;
         LAYER MET3 ;
         RECT  0.0 149.96 180.88 150.52 ;
         LAYER MET3 ;
         RECT  125.12 199.64 682.28 200.2 ;
         LAYER MET3 ;
         RECT  178.48 497.72 682.28 498.28 ;
         LAYER MET3 ;
         RECT  0.0 13.8 276.56 14.36 ;
         LAYER MET3 ;
         RECT  0.0 319.24 682.28 319.8 ;
         LAYER MET3 ;
         RECT  0.0 118.68 122.92 119.24 ;
         LAYER MET4 ;
         RECT  324.76 0.0 325.32 578.32 ;
         LAYER MET4 ;
         RECT  475.64 0.0 476.2 578.32 ;
         LAYER MET4 ;
         RECT  578.68 0.0 579.24 578.32 ;
         LAYER MET4 ;
         RECT  367.08 0.0 367.64 578.32 ;
         LAYER MET4 ;
         RECT  440.68 0.0 441.24 578.32 ;
         LAYER MET4 ;
         RECT  333.96 0.0 334.52 578.32 ;
         LAYER MET3 ;
         RECT  0.0 278.76 682.28 279.32 ;
         LAYER MET3 ;
         RECT  0.0 115.0 122.92 115.56 ;
         LAYER MET4 ;
         RECT  273.24 0.0 273.8 578.32 ;
         LAYER MET4 ;
         RECT  365.24 6.44 365.8 578.32 ;
         LAYER MET4 ;
         RECT  260.36 13.8 260.92 578.32 ;
         LAYER MET3 ;
         RECT  0.0 449.88 682.28 450.44 ;
         LAYER MET3 ;
         RECT  0.0 527.16 147.76 527.72 ;
         LAYER MET4 ;
         RECT  4.6 0.0 5.16 578.32 ;
         LAYER MET4 ;
         RECT  96.6 0.0 97.16 578.32 ;
         LAYER MET4 ;
         RECT  120.52 0.0 121.08 578.32 ;
         LAYER MET4 ;
         RECT  510.6 0.0 511.16 578.32 ;
         LAYER MET4 ;
         RECT  161.0 0.0 161.56 578.32 ;
         LAYER MET4 ;
         RECT  670.68 0.0 671.24 578.32 ;
         LAYER MET3 ;
         RECT  0.0 155.48 122.92 156.04 ;
         LAYER MET3 ;
         RECT  0.0 306.36 682.28 306.92 ;
         LAYER MET3 ;
         RECT  0.0 431.48 682.28 432.04 ;
         LAYER MET4 ;
         RECT  238.28 0.0 238.84 578.32 ;
         LAYER MET4 ;
         RECT  311.88 26.68 312.44 578.32 ;
         LAYER MET4 ;
         RECT  56.12 0.0 56.68 578.32 ;
         LAYER MET3 ;
         RECT  19.32 91.08 682.28 91.64 ;
         LAYER MET3 ;
         RECT  0.0 230.92 682.28 231.48 ;
         LAYER MET4 ;
         RECT  131.56 0.0 132.12 578.32 ;
         LAYER MET3 ;
         RECT  0.0 420.44 682.28 421.0 ;
         LAYER MET4 ;
         RECT  586.04 0.0 586.6 16.2 ;
         LAYER MET3 ;
         RECT  178.48 126.04 682.28 126.6 ;
         LAYER MET4 ;
         RECT  310.04 15.64 310.6 578.32 ;
         LAYER MET3 ;
         RECT  0.0 521.64 682.28 522.2 ;
         LAYER MET4 ;
         RECT  530.84 0.0 531.4 578.32 ;
         LAYER MET4 ;
         RECT  85.56 0.0 86.12 578.32 ;
         LAYER MET4 ;
         RECT  567.64 0.0 568.2 578.32 ;
         LAYER MET4 ;
         RECT  308.2 0.0 308.76 578.32 ;
         LAYER MET3 ;
         RECT  16.56 70.84 682.28 71.4 ;
         LAYER MET3 ;
         RECT  96.6 80.04 682.28 80.6 ;
         LAYER MET3 ;
         RECT  0.0 532.68 682.28 533.24 ;
         LAYER MET4 ;
         RECT  435.16 0.0 435.72 578.32 ;
         LAYER MET3 ;
         RECT  0.0 199.64 122.92 200.2 ;
         LAYER MET4 ;
         RECT  343.16 26.68 343.72 578.32 ;
         LAYER MET4 ;
         RECT  637.56 0.0 638.12 578.32 ;
         LAYER MET4 ;
         RECT  479.32 0.0 479.88 578.32 ;
         LAYER MET4 ;
         RECT  361.56 0.0 362.12 578.32 ;
         LAYER MET4 ;
         RECT  8.28 0.0 8.84 578.32 ;
         LAYER MET3 ;
         RECT  187.68 85.56 682.28 86.12 ;
         LAYER MET4 ;
         RECT  571.32 0.0 571.88 578.32 ;
         LAYER MET3 ;
         RECT  0.0 512.44 147.76 513.0 ;
         LAYER MET3 ;
         RECT  0.0 471.96 682.28 472.52 ;
         LAYER MET4 ;
         RECT  370.76 45.08 371.32 578.32 ;
         LAYER MET3 ;
         RECT  0.0 245.64 83.36 246.2 ;
         LAYER MET4 ;
         RECT  183.08 6.44 183.64 578.32 ;
         LAYER MET4 ;
         RECT  162.84 0.0 163.4 578.32 ;
         LAYER MET3 ;
         RECT  0.0 153.64 106.36 154.2 ;
         LAYER MET4 ;
         RECT  321.08 0.0 321.64 578.32 ;
         LAYER MET4 ;
         RECT  663.32 0.0 663.88 578.32 ;
         LAYER MET3 ;
         RECT  0.0 541.88 147.76 542.44 ;
         LAYER MET4 ;
         RECT  221.72 26.68 222.28 578.32 ;
         LAYER MET4 ;
         RECT  256.68 0.0 257.24 578.32 ;
         LAYER MET3 ;
         RECT  178.48 398.36 682.28 398.92 ;
         LAYER MET4 ;
         RECT  109.48 0.0 110.04 578.32 ;
         LAYER MET4 ;
         RECT  646.76 26.68 647.32 578.32 ;
         LAYER MET3 ;
         RECT  0.0 501.4 180.88 501.96 ;
         LAYER MET4 ;
         RECT  129.72 0.0 130.28 578.32 ;
         LAYER MET3 ;
         RECT  0.0 317.4 682.28 317.96 ;
         LAYER MET4 ;
         RECT  190.44 0.0 191.0 10.68 ;
         LAYER MET4 ;
         RECT  383.64 0.0 384.2 578.32 ;
         LAYER MET4 ;
         RECT  523.48 45.08 524.04 578.32 ;
         LAYER MET3 ;
         RECT  125.12 120.52 682.28 121.08 ;
         LAYER MET4 ;
         RECT  396.52 0.0 397.08 578.32 ;
         LAYER MET3 ;
         RECT  0.0 8.28 682.28 8.84 ;
         LAYER MET3 ;
         RECT  178.48 225.4 682.28 225.96 ;
         LAYER MET3 ;
         RECT  0.0 197.8 106.36 198.36 ;
         LAYER MET3 ;
         RECT  0.0 227.24 682.28 227.8 ;
         LAYER MET4 ;
         RECT  39.56 0.0 40.12 578.32 ;
         LAYER MET3 ;
         RECT  130.64 133.4 682.28 133.96 ;
         LAYER MET4 ;
         RECT  177.56 11.96 178.12 578.32 ;
         LAYER MET3 ;
         RECT  677.12 78.2 682.28 78.76 ;
         LAYER MET4 ;
         RECT  427.8 0.0 428.36 578.32 ;
         LAYER MET3 ;
         RECT  0.0 505.08 682.28 505.64 ;
         LAYER MET3 ;
         RECT  0.0 435.16 682.28 435.72 ;
         LAYER MET3 ;
         RECT  0.0 269.56 147.76 270.12 ;
         LAYER MET4 ;
         RECT  330.28 0.0 330.84 578.32 ;
         LAYER MET4 ;
         RECT  297.16 0.0 297.72 578.32 ;
         LAYER MET3 ;
         RECT  103.96 271.4 682.28 271.96 ;
         LAYER MET3 ;
         RECT  0.0 573.16 180.88 573.72 ;
         LAYER MET3 ;
         RECT  0.0 23.0 682.28 23.56 ;
         LAYER MET3 ;
         RECT  0.0 299.0 682.28 299.56 ;
         LAYER MET3 ;
         RECT  0.0 4.6 115.56 5.16 ;
         LAYER MET4 ;
         RECT  240.12 0.0 240.68 578.32 ;
         LAYER MET4 ;
         RECT  494.04 0.0 494.6 14.36 ;
         LAYER MET4 ;
         RECT  74.52 0.0 75.08 578.32 ;
         LAYER MET3 ;
         RECT  0.0 352.36 180.88 352.92 ;
         LAYER MET3 ;
         RECT  0.0 129.72 122.92 130.28 ;
         LAYER MET4 ;
         RECT  326.6 0.0 327.16 5.16 ;
         LAYER MET4 ;
         RECT  613.64 0.0 614.2 578.32 ;
         LAYER MET3 ;
         RECT  178.48 282.44 682.28 283.0 ;
         LAYER MET4 ;
         RECT  508.76 0.0 509.32 578.32 ;
         LAYER MET3 ;
         RECT  0.0 538.2 180.88 538.76 ;
         LAYER MET3 ;
         RECT  151.8 92.92 682.28 93.48 ;
         LAYER MET4 ;
         RECT  115.0 0.0 115.56 578.32 ;
         LAYER MET3 ;
         RECT  178.48 57.96 682.28 58.52 ;
         LAYER MET4 ;
         RECT  146.28 0.0 146.84 578.32 ;
         LAYER MET4 ;
         RECT  81.88 0.0 82.44 578.32 ;
         LAYER MET3 ;
         RECT  178.48 425.96 682.28 426.52 ;
         LAYER MET4 ;
         RECT  540.04 0.0 540.6 578.32 ;
         LAYER MET3 ;
         RECT  0.0 343.16 682.28 343.72 ;
         LAYER MET4 ;
         RECT  67.16 0.0 67.72 578.32 ;
         LAYER MET4 ;
         RECT  446.2 0.0 446.76 578.32 ;
         LAYER MET4 ;
         RECT  133.4 0.0 133.96 578.32 ;
         LAYER MET4 ;
         RECT  560.28 0.0 560.84 578.32 ;
         LAYER MET3 ;
         RECT  0.0 392.84 682.28 393.4 ;
         LAYER MET3 ;
         RECT  0.0 35.88 119.24 36.44 ;
         LAYER MET4 ;
         RECT  514.28 0.0 514.84 578.32 ;
         LAYER MET4 ;
         RECT  2.76 0.0 3.32 578.32 ;
         LAYER MET4 ;
         RECT  400.2 0.0 400.76 578.32 ;
         LAYER MET3 ;
         RECT  0.0 221.72 122.92 222.28 ;
         LAYER MET3 ;
         RECT  0.0 236.44 180.88 237.0 ;
         LAYER MET4 ;
         RECT  319.24 0.0 319.8 578.32 ;
         LAYER MET3 ;
         RECT  0.0 238.28 83.36 238.84 ;
         LAYER MET3 ;
         RECT  0.0 253.0 682.28 253.56 ;
         LAYER MET4 ;
         RECT  124.2 0.0 124.76 578.32 ;
         LAYER MET4 ;
         RECT  194.12 0.0 194.68 5.16 ;
         LAYER MET3 ;
         RECT  96.6 61.64 682.28 62.2 ;
         LAYER MET3 ;
         RECT  0.0 488.52 682.28 489.08 ;
         LAYER MET3 ;
         RECT  178.48 527.16 682.28 527.72 ;
         LAYER MET4 ;
         RECT  253.0 0.0 253.56 578.32 ;
         LAYER MET3 ;
         RECT  0.0 184.92 682.28 185.48 ;
         LAYER MET3 ;
         RECT  0.0 567.64 682.28 568.2 ;
         LAYER MET4 ;
         RECT  72.68 0.0 73.24 578.32 ;
         LAYER MET4 ;
         RECT  276.92 15.64 277.48 578.32 ;
         LAYER MET3 ;
         RECT  0.0 374.44 682.28 375.0 ;
         LAYER MET4 ;
         RECT  556.6 0.0 557.16 578.32 ;
         LAYER MET4 ;
         RECT  576.84 0.0 577.4 578.32 ;
         LAYER MET4 ;
         RECT  517.96 0.0 518.52 578.32 ;
         LAYER MET4 ;
         RECT  494.04 26.68 494.6 578.32 ;
         LAYER MET3 ;
         RECT  0.0 207.0 122.92 207.56 ;
         LAYER MET3 ;
         RECT  0.0 376.28 682.28 376.84 ;
         LAYER MET4 ;
         RECT  519.8 0.0 520.36 578.32 ;
         LAYER MET4 ;
         RECT  563.96 0.0 564.52 578.32 ;
         LAYER MET3 ;
         RECT  0.0 400.2 682.28 400.76 ;
         LAYER MET3 ;
         RECT  100.28 238.28 682.28 238.84 ;
         LAYER MET3 ;
         RECT  0.0 302.68 682.28 303.24 ;
         LAYER MET3 ;
         RECT  0.0 543.72 682.28 544.28 ;
         LAYER MET4 ;
         RECT  113.16 0.0 113.72 578.32 ;
         LAYER MET4 ;
         RECT  11.96 0.0 12.52 578.32 ;
         LAYER MET3 ;
         RECT  0.0 460.92 682.28 461.48 ;
         LAYER MET4 ;
         RECT  59.8 0.0 60.36 578.32 ;
         LAYER MET4 ;
         RECT  525.32 0.0 525.88 10.68 ;
         LAYER MET3 ;
         RECT  0.0 517.96 682.28 518.52 ;
         LAYER MET3 ;
         RECT  0.0 208.84 122.92 209.4 ;
         LAYER MET3 ;
         RECT  0.0 168.36 106.36 168.92 ;
         LAYER MET4 ;
         RECT  219.88 0.0 220.44 578.32 ;
         LAYER MET4 ;
         RECT  168.36 0.0 168.92 578.32 ;
         LAYER MET3 ;
         RECT  0.0 361.56 682.28 362.12 ;
         LAYER MET3 ;
         RECT  0.0 523.48 180.88 524.04 ;
         LAYER MET3 ;
         RECT  0.0 21.16 682.28 21.72 ;
         LAYER MET4 ;
         RECT  385.48 0.0 386.04 578.32 ;
         LAYER MET4 ;
         RECT  69.0 0.0 69.56 578.32 ;
         LAYER MET3 ;
         RECT  0.0 186.76 180.88 187.32 ;
         LAYER MET4 ;
         RECT  455.4 0.0 455.96 578.32 ;
         LAYER MET4 ;
         RECT  181.24 0.0 181.8 578.32 ;
         LAYER MET3 ;
         RECT  125.12 113.16 682.28 113.72 ;
         LAYER MET3 ;
         RECT  0.0 120.52 7.0 121.08 ;
         LAYER MET3 ;
         RECT  0.0 232.76 682.28 233.32 ;
         LAYER MET3 ;
         RECT  0.0 219.88 122.92 220.44 ;
         LAYER MET4 ;
         RECT  212.52 0.0 213.08 578.32 ;
         LAYER MET4 ;
         RECT  665.16 0.0 665.72 578.32 ;
         LAYER MET4 ;
         RECT  376.28 0.0 376.84 5.16 ;
         LAYER MET3 ;
         RECT  0.0 483.0 682.28 483.56 ;
         LAYER MET4 ;
         RECT  243.8 13.8 244.36 578.32 ;
         LAYER MET4 ;
         RECT  394.68 0.0 395.24 578.32 ;
         LAYER MET3 ;
         RECT  101.2 245.64 682.28 246.2 ;
         LAYER MET4 ;
         RECT  589.72 0.0 590.28 578.32 ;
         LAYER MET3 ;
         RECT  0.0 214.36 122.92 214.92 ;
         LAYER MET4 ;
         RECT  223.56 0.0 224.12 578.32 ;
         LAYER MET3 ;
         RECT  0.0 563.96 682.28 564.52 ;
         LAYER MET3 ;
         RECT  177.56 76.36 682.28 76.92 ;
         LAYER MET4 ;
         RECT  672.52 0.0 673.08 578.32 ;
         LAYER MET4 ;
         RECT  282.44 26.68 283.0 578.32 ;
         LAYER MET3 ;
         RECT  427.8 2.76 682.28 3.32 ;
         LAYER MET4 ;
         RECT  267.72 0.0 268.28 578.32 ;
         LAYER MET3 ;
         RECT  0.0 111.32 106.36 111.88 ;
         LAYER MET4 ;
         RECT  547.4 0.0 547.96 578.32 ;
         LAYER MET4 ;
         RECT  87.4 0.0 87.96 578.32 ;
         LAYER MET4 ;
         RECT  354.2 0.0 354.76 578.32 ;
         LAYER MET3 ;
         RECT  39.56 32.2 682.28 32.76 ;
         LAYER MET4 ;
         RECT  57.96 0.0 58.52 578.32 ;
         LAYER MET3 ;
         RECT  0.0 378.12 682.28 378.68 ;
         LAYER MET4 ;
         RECT  230.92 0.0 231.48 578.32 ;
         LAYER MET4 ;
         RECT  245.64 0.0 246.2 578.32 ;
         LAYER MET4 ;
         RECT  78.2 0.0 78.76 578.32 ;
         LAYER MET4 ;
         RECT  405.72 0.0 406.28 578.32 ;
         LAYER MET4 ;
         RECT  549.24 0.0 549.8 578.32 ;
         LAYER MET3 ;
         RECT  0.0 468.28 682.28 468.84 ;
         LAYER MET3 ;
         RECT  0.0 103.96 7.0 104.52 ;
         LAYER MET4 ;
         RECT  593.4 0.0 593.96 578.32 ;
         LAYER MET3 ;
         RECT  0.0 370.76 682.28 371.32 ;
         LAYER MET3 ;
         RECT  0.0 470.12 147.76 470.68 ;
         LAYER MET3 ;
         RECT  0.0 348.68 682.28 349.24 ;
         LAYER MET3 ;
         RECT  0.0 499.56 682.28 500.12 ;
         LAYER MET3 ;
         RECT  0.0 291.64 682.28 292.2 ;
         LAYER MET3 ;
         RECT  0.0 385.48 682.28 386.04 ;
         LAYER MET4 ;
         RECT  251.16 26.68 251.72 578.32 ;
         LAYER MET4 ;
         RECT  503.24 0.0 503.8 578.32 ;
         LAYER MET3 ;
         RECT  0.0 240.12 147.76 240.68 ;
         LAYER MET3 ;
         RECT  132.48 19.32 682.28 19.88 ;
         LAYER MET3 ;
         RECT  19.32 124.2 682.28 124.76 ;
         LAYER MET3 ;
         RECT  178.48 354.2 682.28 354.76 ;
         LAYER MET4 ;
         RECT  306.36 0.0 306.92 578.32 ;
         LAYER MET4 ;
         RECT  216.2 6.44 216.76 578.32 ;
         LAYER MET3 ;
         RECT  178.48 512.44 682.28 513.0 ;
         LAYER MET4 ;
         RECT  580.52 0.0 581.08 578.32 ;
         LAYER MET3 ;
         RECT  0.0 273.24 180.88 273.8 ;
         LAYER MET4 ;
         RECT  241.96 0.0 242.52 578.32 ;
         LAYER MET4 ;
         RECT  363.4 0.0 363.96 578.32 ;
         LAYER MET4 ;
         RECT  499.56 0.0 500.12 578.32 ;
         LAYER MET4 ;
         RECT  444.36 0.0 444.92 578.32 ;
         LAYER MET4 ;
         RECT  94.76 0.0 95.32 578.32 ;
         LAYER MET3 ;
         RECT  178.48 413.08 682.28 413.64 ;
         LAYER MET4 ;
         RECT  630.2 0.0 630.76 578.32 ;
         LAYER MET4 ;
         RECT  10.12 0.0 10.68 578.32 ;
         LAYER MET4 ;
         RECT  122.36 0.0 122.92 578.32 ;
         LAYER MET4 ;
         RECT  70.84 0.0 71.4 578.32 ;
         LAYER MET4 ;
         RECT  48.76 0.0 49.32 578.32 ;
         LAYER MET4 ;
         RECT  262.2 0.0 262.76 578.32 ;
         LAYER MET4 ;
         RECT  387.32 0.0 387.88 578.32 ;
         LAYER MET3 ;
         RECT  0.0 464.6 682.28 465.16 ;
         LAYER MET4 ;
         RECT  254.84 0.0 255.4 578.32 ;
         LAYER MET3 ;
         RECT  0.0 324.76 682.28 325.32 ;
         LAYER MET3 ;
         RECT  132.48 161.0 682.28 161.56 ;
         LAYER MET3 ;
         RECT  89.24 241.96 682.28 242.52 ;
         LAYER MET3 ;
         RECT  0.0 105.8 682.28 106.36 ;
         LAYER MET3 ;
         RECT  178.48 326.6 682.28 327.16 ;
         LAYER MET4 ;
         RECT  648.6 0.0 649.16 578.32 ;
         LAYER MET3 ;
         RECT  16.56 103.96 682.28 104.52 ;
         LAYER MET3 ;
         RECT  0.0 497.72 147.76 498.28 ;
         LAYER MET4 ;
         RECT  63.48 0.0 64.04 578.32 ;
         LAYER MET3 ;
         RECT  178.48 183.08 682.28 183.64 ;
         LAYER MET4 ;
         RECT  61.64 0.0 62.2 578.32 ;
         LAYER MET3 ;
         RECT  0.0 161.0 122.92 161.56 ;
         LAYER MET3 ;
         RECT  0.0 356.04 682.28 356.6 ;
         LAYER MET3 ;
         RECT  0.0 413.08 147.76 413.64 ;
         LAYER MET3 ;
         RECT  0.0 300.84 180.88 301.4 ;
         LAYER MET3 ;
         RECT  0.0 19.32 119.24 19.88 ;
         LAYER MET3 ;
         RECT  136.16 205.16 682.28 205.72 ;
         LAYER MET4 ;
         RECT  207.0 0.0 207.56 578.32 ;
         LAYER MET4 ;
         RECT  348.68 6.44 349.24 578.32 ;
         LAYER MET4 ;
         RECT  532.68 0.0 533.24 578.32 ;
         LAYER MET4 ;
         RECT  650.44 0.0 651.0 578.32 ;
         LAYER MET3 ;
         RECT  0.0 262.2 682.28 262.76 ;
         LAYER MET4 ;
         RECT  105.8 0.0 106.36 578.32 ;
         LAYER MET4 ;
         RECT  425.96 19.32 426.52 578.32 ;
         LAYER MET3 ;
         RECT  0.0 394.68 180.88 395.24 ;
         LAYER MET4 ;
         RECT  409.4 11.96 409.96 578.32 ;
         LAYER MET3 ;
         RECT  0.0 177.56 122.92 178.12 ;
         LAYER MET3 ;
         RECT  0.0 39.56 22.64 40.12 ;
         LAYER MET4 ;
         RECT  431.48 45.08 432.04 578.32 ;
         LAYER MET4 ;
         RECT  15.64 0.0 16.2 578.32 ;
         LAYER MET3 ;
         RECT  0.0 256.68 682.28 257.24 ;
         LAYER MET4 ;
         RECT  293.48 11.96 294.04 578.32 ;
         LAYER MET3 ;
         RECT  0.0 183.08 106.36 183.64 ;
         LAYER MET4 ;
         RECT  24.84 0.0 25.4 578.32 ;
         LAYER MET3 ;
         RECT  0.0 34.04 22.64 34.6 ;
         LAYER MET4 ;
         RECT  151.8 0.0 152.36 578.32 ;
         LAYER MET3 ;
         RECT  0.0 422.28 682.28 422.84 ;
         LAYER MET3 ;
         RECT  132.48 35.88 682.28 36.44 ;
         LAYER MET3 ;
         RECT  0.0 335.8 682.28 336.36 ;
         LAYER MET3 ;
         RECT  0.0 407.56 682.28 408.12 ;
         LAYER MET3 ;
         RECT  0.0 529.0 682.28 529.56 ;
         LAYER MET4 ;
         RECT  289.8 0.0 290.36 578.32 ;
         LAYER MET4 ;
         RECT  135.24 0.0 135.8 578.32 ;
         LAYER MET4 ;
         RECT  527.16 0.0 527.72 578.32 ;
         LAYER MET4 ;
         RECT  529.0 0.0 529.56 578.32 ;
         LAYER MET3 ;
         RECT  0.0 381.8 682.28 382.36 ;
         LAYER MET3 ;
         RECT  0.0 558.44 180.88 559.0 ;
         LAYER MET4 ;
         RECT  538.2 0.0 538.76 578.32 ;
         LAYER MET3 ;
         RECT  427.8 6.44 682.28 7.0 ;
         LAYER MET3 ;
         RECT  0.0 286.12 180.88 286.68 ;
         LAYER MET3 ;
         RECT  0.0 519.8 682.28 520.36 ;
         LAYER MET3 ;
         RECT  0.0 495.88 682.28 496.44 ;
         LAYER MET4 ;
         RECT  611.8 0.0 612.36 578.32 ;
         LAYER MET3 ;
         RECT  0.0 54.28 682.28 54.84 ;
         LAYER MET4 ;
         RECT  280.6 0.0 281.16 578.32 ;
         LAYER MET3 ;
         RECT  125.12 135.24 682.28 135.8 ;
         LAYER MET4 ;
         RECT  300.84 0.0 301.4 578.32 ;
         LAYER MET4 ;
         RECT  654.12 0.0 654.68 578.32 ;
         LAYER MET3 ;
         RECT  0.0 59.8 191.92 60.36 ;
         LAYER MET3 ;
         RECT  103.04 264.04 682.28 264.6 ;
         LAYER MET3 ;
         RECT  19.32 74.52 682.28 75.08 ;
         LAYER MET4 ;
         RECT  598.92 0.0 599.48 578.32 ;
         LAYER MET4 ;
         RECT  429.64 0.0 430.2 578.32 ;
         LAYER MET4 ;
         RECT  118.68 0.0 119.24 578.32 ;
         LAYER MET3 ;
         RECT  125.12 212.52 682.28 213.08 ;
         LAYER MET3 ;
         RECT  0.0 102.12 682.28 102.68 ;
         LAYER MET4 ;
         RECT  413.08 0.0 413.64 578.32 ;
         LAYER MET4 ;
         RECT  332.12 0.0 332.68 578.32 ;
         LAYER MET3 ;
         RECT  0.0 188.6 682.28 189.16 ;
         LAYER MET3 ;
         RECT  0.0 571.32 179.04 571.88 ;
         LAYER MET4 ;
         RECT  299.0 6.44 299.56 578.32 ;
         LAYER MET4 ;
         RECT  225.4 0.0 225.96 578.32 ;
         LAYER MET3 ;
         RECT  0.0 560.28 682.28 560.84 ;
         LAYER MET4 ;
         RECT  409.4 0.0 409.96 5.16 ;
         LAYER MET3 ;
         RECT  0.0 534.52 682.28 535.08 ;
         LAYER MET4 ;
         RECT  173.88 0.0 174.44 578.32 ;
         LAYER MET3 ;
         RECT  0.0 126.04 106.36 126.6 ;
         LAYER MET4 ;
         RECT  275.08 0.0 275.64 578.32 ;
         LAYER MET4 ;
         RECT  641.24 0.0 641.8 578.32 ;
         LAYER MET3 ;
         RECT  0.0 275.08 682.28 275.64 ;
         LAYER MET3 ;
         RECT  0.0 330.28 180.88 330.84 ;
         LAYER MET3 ;
         RECT  0.0 446.2 682.28 446.76 ;
         LAYER MET4 ;
         RECT  284.28 0.0 284.84 578.32 ;
         LAYER MET3 ;
         RECT  0.0 223.56 682.28 224.12 ;
         LAYER MET4 ;
         RECT  403.88 26.68 404.44 578.32 ;
         LAYER MET3 ;
         RECT  495.88 15.64 682.28 16.2 ;
         LAYER MET4 ;
         RECT  632.04 0.0 632.6 578.32 ;
         LAYER MET4 ;
         RECT  137.08 0.0 137.64 578.32 ;
         LAYER MET3 ;
         RECT  0.0 565.8 180.88 566.36 ;
         LAYER MET4 ;
         RECT  142.6 0.0 143.16 578.32 ;
         LAYER MET4 ;
         RECT  575.0 0.0 575.56 578.32 ;
         LAYER MET3 ;
         RECT  0.0 70.84 7.0 71.4 ;
         LAYER MET4 ;
         RECT  407.56 0.0 408.12 578.32 ;
         LAYER MET3 ;
         RECT  0.0 459.08 180.88 459.64 ;
         LAYER MET4 ;
         RECT  389.16 0.0 389.72 578.32 ;
         LAYER MET3 ;
         RECT  132.48 52.44 682.28 53.0 ;
         LAYER MET3 ;
         RECT  0.0 350.52 682.28 351.08 ;
         LAYER MET3 ;
         RECT  96.6 45.08 682.28 45.64 ;
         LAYER MET3 ;
         RECT  0.0 284.28 682.28 284.84 ;
         LAYER MET4 ;
         RECT  310.04 0.0 310.6 5.16 ;
         LAYER MET3 ;
         RECT  0.0 72.68 682.28 73.24 ;
         LAYER MET4 ;
         RECT  619.16 0.0 619.72 578.32 ;
         LAYER MET3 ;
         RECT  0.0 368.92 147.76 369.48 ;
         LAYER MET3 ;
         RECT  0.0 0.92 119.24 1.48 ;
         LAYER MET4 ;
         RECT  89.24 0.0 89.8 578.32 ;
         LAYER MET3 ;
         RECT  420.44 0.92 682.28 1.48 ;
         LAYER MET3 ;
         RECT  0.0 536.36 682.28 536.92 ;
         LAYER MET3 ;
         RECT  0.0 46.92 682.28 47.48 ;
         LAYER MET4 ;
         RECT  606.28 0.0 606.84 578.32 ;
         LAYER MET3 ;
         RECT  416.76 4.6 682.28 5.16 ;
         LAYER MET4 ;
         RECT  92.92 0.0 93.48 578.32 ;
         LAYER MET3 ;
         RECT  0.0 304.52 682.28 305.08 ;
         LAYER MET4 ;
         RECT  536.36 0.0 536.92 578.32 ;
         LAYER MET3 ;
         RECT  178.48 297.16 682.28 297.72 ;
         LAYER MET3 ;
         RECT  650.44 59.8 682.28 60.36 ;
         LAYER MET3 ;
         RECT  0.0 438.84 682.28 439.4 ;
         LAYER MET4 ;
         RECT  172.04 0.0 172.6 578.32 ;
         LAYER MET4 ;
         RECT  103.96 0.0 104.52 578.32 ;
         LAYER MET4 ;
         RECT  483.0 0.0 483.56 578.32 ;
         LAYER MET4 ;
         RECT  343.16 0.0 343.72 5.16 ;
         LAYER MET3 ;
         RECT  0.0 56.12 682.28 56.68 ;
         LAYER MET3 ;
         RECT  0.0 181.24 682.28 181.8 ;
         LAYER MET3 ;
         RECT  0.0 367.08 682.28 367.64 ;
         LAYER MET4 ;
         RECT  175.72 0.0 176.28 578.32 ;
         LAYER MET4 ;
         RECT  552.92 0.0 553.48 578.32 ;
         LAYER MET3 ;
         RECT  0.0 552.92 180.88 553.48 ;
         LAYER MET3 ;
         RECT  0.0 146.28 682.28 146.84 ;
         LAYER MET3 ;
         RECT  0.0 89.24 682.28 89.8 ;
         LAYER MET3 ;
         RECT  0.0 289.8 682.28 290.36 ;
         LAYER MET3 ;
         RECT  0.0 251.16 180.88 251.72 ;
         LAYER MET4 ;
         RECT  628.36 0.0 628.92 578.32 ;
         LAYER MET3 ;
         RECT  16.56 87.4 682.28 87.96 ;
         LAYER MET3 ;
         RECT  0.0 142.6 180.88 143.16 ;
         LAYER MET4 ;
         RECT  17.48 0.0 18.04 578.32 ;
         LAYER MET3 ;
         RECT  0.0 216.2 682.28 216.76 ;
         LAYER MET4 ;
         RECT  341.32 0.0 341.88 578.32 ;
         LAYER MET3 ;
         RECT  178.48 269.56 682.28 270.12 ;
         LAYER MET3 ;
         RECT  0.0 144.44 682.28 145.0 ;
         LAYER MET4 ;
         RECT  45.08 0.0 45.64 578.32 ;
         LAYER MET4 ;
         RECT  486.68 0.0 487.24 578.32 ;
         LAYER MET4 ;
         RECT  569.48 0.0 570.04 578.32 ;
         LAYER MET4 ;
         RECT  609.96 0.0 610.52 578.32 ;
         LAYER MET4 ;
         RECT  227.24 0.0 227.8 5.16 ;
         LAYER MET3 ;
         RECT  0.0 425.96 147.76 426.52 ;
         LAYER MET4 ;
         RECT  30.36 0.0 30.92 578.32 ;
         LAYER MET4 ;
         RECT  203.32 0.0 203.88 578.32 ;
         LAYER MET4 ;
         RECT  286.12 0.0 286.68 578.32 ;
         LAYER MET4 ;
         RECT  157.32 0.0 157.88 578.32 ;
         LAYER MET4 ;
         RECT  608.12 0.0 608.68 578.32 ;
         LAYER MET3 ;
         RECT  0.0 276.92 86.12 277.48 ;
         LAYER MET3 ;
         RECT  178.48 484.84 682.28 485.4 ;
         LAYER MET4 ;
         RECT  243.8 0.0 244.36 5.16 ;
         LAYER MET3 ;
         RECT  0.0 148.12 682.28 148.68 ;
         LAYER MET3 ;
         RECT  0.0 540.04 682.28 540.6 ;
         LAYER MET4 ;
         RECT  595.24 0.0 595.8 578.32 ;
         LAYER MET3 ;
         RECT  0.0 172.04 122.92 172.6 ;
         LAYER MET4 ;
         RECT  37.72 33.12 38.28 578.32 ;
         LAYER MET3 ;
         RECT  0.0 554.76 682.28 555.32 ;
         LAYER MET4 ;
         RECT  551.08 0.0 551.64 578.32 ;
         LAYER MET4 ;
         RECT  652.28 0.0 652.84 578.32 ;
         LAYER MET3 ;
         RECT  178.48 210.68 682.28 211.24 ;
         LAYER MET4 ;
         RECT  420.44 0.0 421.0 578.32 ;
         LAYER MET3 ;
         RECT  0.0 243.8 180.88 244.36 ;
         LAYER MET3 ;
         RECT  0.0 451.72 180.88 452.28 ;
         LAYER MET3 ;
         RECT  0.0 122.36 122.92 122.92 ;
         LAYER MET4 ;
         RECT  411.24 0.0 411.8 578.32 ;
         LAYER MET4 ;
         RECT  28.52 0.0 29.08 578.32 ;
         LAYER MET4 ;
         RECT  247.48 0.0 248.04 578.32 ;
         LAYER MET3 ;
         RECT  0.0 190.44 682.28 191.0 ;
         LAYER MET3 ;
         RECT  0.0 11.96 210.32 12.52 ;
         LAYER MET4 ;
         RECT  127.88 0.0 128.44 578.32 ;
         LAYER MET4 ;
         RECT  227.24 11.96 227.8 578.32 ;
         LAYER MET3 ;
         RECT  0.0 137.08 7.0 137.64 ;
         LAYER MET4 ;
         RECT  265.88 6.44 266.44 578.32 ;
         LAYER MET3 ;
         RECT  0.0 78.2 191.92 78.76 ;
         LAYER MET3 ;
         RECT  0.0 494.04 180.88 494.6 ;
         LAYER MET3 ;
         RECT  526.24 11.96 682.28 12.52 ;
         LAYER MET3 ;
         RECT  19.32 83.72 682.28 84.28 ;
         LAYER MET3 ;
         RECT  0.0 131.56 682.28 132.12 ;
         LAYER MET3 ;
         RECT  0.0 332.12 682.28 332.68 ;
         LAYER MET4 ;
         RECT  140.76 0.0 141.32 578.32 ;
         LAYER MET4 ;
         RECT  543.72 0.0 544.28 578.32 ;
         LAYER MET3 ;
         RECT  0.0 195.96 682.28 196.52 ;
         LAYER MET3 ;
         RECT  0.0 549.24 682.28 549.8 ;
         LAYER MET3 ;
         RECT  0.0 96.6 93.48 97.16 ;
         LAYER MET4 ;
         RECT  490.36 0.0 490.92 578.32 ;
         LAYER MET4 ;
         RECT  374.44 0.0 375.0 578.32 ;
         LAYER MET4 ;
         RECT  194.12 11.96 194.68 578.32 ;
         LAYER MET3 ;
         RECT  125.12 177.56 682.28 178.12 ;
         LAYER MET3 ;
         RECT  0.0 69.0 119.24 69.56 ;
         LAYER MET3 ;
         RECT  0.0 455.4 147.76 455.96 ;
         LAYER MET3 ;
         RECT  125.12 219.88 682.28 220.44 ;
         LAYER MET4 ;
         RECT  391.0 0.0 391.56 578.32 ;
         LAYER MET3 ;
         RECT  96.6 96.6 682.28 97.16 ;
         LAYER MET4 ;
         RECT  438.84 0.0 439.4 578.32 ;
         LAYER MET3 ;
         RECT  178.48 440.68 682.28 441.24 ;
         LAYER MET3 ;
         RECT  0.0 525.32 682.28 525.88 ;
         LAYER MET3 ;
         RECT  178.48 311.88 682.28 312.44 ;
         LAYER MET4 ;
         RECT  376.28 15.64 376.84 578.32 ;
         LAYER MET3 ;
         RECT  0.0 135.24 122.92 135.8 ;
         LAYER MET4 ;
         RECT  190.44 26.68 191.0 578.32 ;
         LAYER MET4 ;
         RECT  26.68 0.0 27.24 578.32 ;
         LAYER MET4 ;
         RECT  488.52 0.0 489.08 578.32 ;
         LAYER MET3 ;
         RECT  125.12 127.88 682.28 128.44 ;
         LAYER MET3 ;
         RECT  0.0 287.96 682.28 288.52 ;
         LAYER MET4 ;
         RECT  221.72 0.0 222.28 10.68 ;
         LAYER MET3 ;
         RECT  0.0 313.72 682.28 314.28 ;
         LAYER MET3 ;
         RECT  0.0 556.6 147.76 557.16 ;
         LAYER MET4 ;
         RECT  210.68 0.0 211.24 5.16 ;
         LAYER MET3 ;
         RECT  0.0 530.84 180.88 531.4 ;
         LAYER MET4 ;
         RECT  484.84 0.0 485.4 578.32 ;
         LAYER MET3 ;
         RECT  0.0 326.6 147.76 327.16 ;
         LAYER MET4 ;
         RECT  451.72 0.0 452.28 578.32 ;
         LAYER MET3 ;
         RECT  0.0 322.92 180.88 323.48 ;
         LAYER MET3 ;
         RECT  0.0 490.36 682.28 490.92 ;
         LAYER MET3 ;
         RECT  0.0 15.64 342.8 16.2 ;
         LAYER MET3 ;
         RECT  0.0 473.8 180.88 474.36 ;
         LAYER MET4 ;
         RECT  626.52 0.0 627.08 578.32 ;
         LAYER MET4 ;
         RECT  359.72 13.8 360.28 578.32 ;
         LAYER MET3 ;
         RECT  0.0 477.48 682.28 478.04 ;
         LAYER MET3 ;
         RECT  0.0 508.76 180.88 509.32 ;
         LAYER MET4 ;
         RECT  591.56 0.0 592.12 578.32 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER MET3 ;
         RECT  0.0 309.12 182.72 309.68 ;
         LAYER MET3 ;
         RECT  81.88 29.44 682.28 30.0 ;
         LAYER MET3 ;
         RECT  0.0 97.52 682.28 98.08 ;
         LAYER MET3 ;
         RECT  0.0 390.08 147.76 390.64 ;
         LAYER MET4 ;
         RECT  553.84 45.08 554.4 578.32 ;
         LAYER MET3 ;
         RECT  678.96 408.48 682.28 409.04 ;
         LAYER MET3 ;
         RECT  50.6 38.64 682.28 39.2 ;
         LAYER MET3 ;
         RECT  0.0 169.28 122.92 169.84 ;
         LAYER MET3 ;
         RECT  0.0 448.96 147.76 449.52 ;
         LAYER MET4 ;
         RECT  634.8 0.0 635.36 578.32 ;
         LAYER MET3 ;
         RECT  678.96 566.72 682.28 567.28 ;
         LAYER MET4 ;
         RECT  671.6 0.0 672.16 578.32 ;
         LAYER MET4 ;
         RECT  11.04 0.0 11.6 578.32 ;
         LAYER MET3 ;
         RECT  187.68 84.64 682.28 85.2 ;
         LAYER MET3 ;
         RECT  0.0 9.2 119.24 9.76 ;
         LAYER MET3 ;
         RECT  678.96 494.96 682.28 495.52 ;
         LAYER MET3 ;
         RECT  678.96 121.44 682.28 122.0 ;
         LAYER MET4 ;
         RECT  36.8 33.12 37.36 578.32 ;
         LAYER MET4 ;
         RECT  241.04 0.0 241.6 578.32 ;
         LAYER MET4 ;
         RECT  310.96 15.64 311.52 578.32 ;
         LAYER MET4 ;
         RECT  572.24 0.0 572.8 578.32 ;
         LAYER MET4 ;
         RECT  228.16 0.0 228.72 5.16 ;
         LAYER MET3 ;
         RECT  678.96 452.64 682.28 453.2 ;
         LAYER MET3 ;
         RECT  0.0 64.4 682.28 64.96 ;
         LAYER MET4 ;
         RECT  375.36 0.0 375.92 578.32 ;
         LAYER MET3 ;
         RECT  0.0 537.28 182.72 537.84 ;
         LAYER MET3 ;
         RECT  678.96 114.08 682.28 114.64 ;
         LAYER MET3 ;
         RECT  678.96 574.08 682.28 574.64 ;
         LAYER MET4 ;
         RECT  555.68 0.0 556.24 12.52 ;
         LAYER MET3 ;
         RECT  0.0 279.68 182.72 280.24 ;
         LAYER MET3 ;
         RECT  0.0 292.56 682.28 293.12 ;
         LAYER MET3 ;
         RECT  0.0 228.16 78.76 228.72 ;
         LAYER MET3 ;
         RECT  0.0 329.36 182.72 329.92 ;
         LAYER MET4 ;
         RECT  568.56 0.0 569.12 578.32 ;
         LAYER MET3 ;
         RECT  0.0 235.52 682.28 236.08 ;
         LAYER MET4 ;
         RECT  134.32 6.44 134.88 578.32 ;
         LAYER MET4 ;
         RECT  130.64 0.0 131.2 578.32 ;
         LAYER MET4 ;
         RECT  496.8 0.0 497.36 578.32 ;
         LAYER MET3 ;
         RECT  678.96 472.88 682.28 473.44 ;
         LAYER MET4 ;
         RECT  90.16 0.0 90.72 578.32 ;
         LAYER MET3 ;
         RECT  0.0 44.16 25.4 44.72 ;
         LAYER MET4 ;
         RECT  9.2 0.0 9.76 578.32 ;
         LAYER MET4 ;
         RECT  29.44 0.0 30.0 578.32 ;
         LAYER MET3 ;
         RECT  129.72 125.12 682.28 125.68 ;
         LAYER MET3 ;
         RECT  178.48 132.48 682.28 133.04 ;
         LAYER MET3 ;
         RECT  178.48 233.68 682.28 234.24 ;
         LAYER MET4 ;
         RECT  112.24 0.0 112.8 578.32 ;
         LAYER MET4 ;
         RECT  417.68 0.0 418.24 578.32 ;
         LAYER MET4 ;
         RECT  552.0 0.0 552.56 578.32 ;
         LAYER MET4 ;
         RECT  138.0 0.0 138.56 578.32 ;
         LAYER MET3 ;
         RECT  89.24 266.8 682.28 267.36 ;
         LAYER MET3 ;
         RECT  0.0 283.36 682.28 283.92 ;
         LAYER MET4 ;
         RECT  432.4 45.08 432.96 578.32 ;
         LAYER MET4 ;
         RECT  336.72 0.0 337.28 578.32 ;
         LAYER MET4 ;
         RECT  393.76 0.0 394.32 5.16 ;
         LAYER MET3 ;
         RECT  0.0 307.28 682.28 307.84 ;
         LAYER MET4 ;
         RECT  590.64 0.0 591.2 578.32 ;
         LAYER MET4 ;
         RECT  581.44 0.0 582.0 578.32 ;
         LAYER MET4 ;
         RECT  384.56 0.0 385.12 578.32 ;
         LAYER MET4 ;
         RECT  364.32 6.44 364.88 578.32 ;
         LAYER MET3 ;
         RECT  0.0 233.68 86.12 234.24 ;
         LAYER MET3 ;
         RECT  0.0 217.12 682.28 217.68 ;
         LAYER MET3 ;
         RECT  0.0 322.0 182.72 322.56 ;
         LAYER MET3 ;
         RECT  678.96 250.24 682.28 250.8 ;
         LAYER MET4 ;
         RECT  1.84 0.0 2.4 84.28 ;
         LAYER MET3 ;
         RECT  0.0 496.8 682.28 497.36 ;
         LAYER MET4 ;
         RECT  16.56 0.0 17.12 578.32 ;
         LAYER MET4 ;
         RECT  235.52 0.0 236.08 578.32 ;
         LAYER MET3 ;
         RECT  0.0 507.84 682.28 508.4 ;
         LAYER MET4 ;
         RECT  34.96 0.0 35.52 578.32 ;
         LAYER MET4 ;
         RECT  408.48 0.0 409.04 578.32 ;
         LAYER MET3 ;
         RECT  0.0 193.2 182.72 193.76 ;
         LAYER MET3 ;
         RECT  0.0 517.04 182.72 517.6 ;
         LAYER MET4 ;
         RECT  136.16 0.0 136.72 578.32 ;
         LAYER MET3 ;
         RECT  0.0 160.08 682.28 160.64 ;
         LAYER MET3 ;
         RECT  0.0 207.92 122.92 208.48 ;
         LAYER MET3 ;
         RECT  0.0 467.36 682.28 467.92 ;
         LAYER MET3 ;
         RECT  0.0 471.04 682.28 471.6 ;
         LAYER MET3 ;
         RECT  0.0 386.4 182.72 386.96 ;
         LAYER MET4 ;
         RECT  231.84 6.44 232.4 578.32 ;
         LAYER MET4 ;
         RECT  428.72 0.0 429.28 578.32 ;
         LAYER MET4 ;
         RECT  588.8 0.0 589.36 578.32 ;
         LAYER MET3 ;
         RECT  0.0 277.84 682.28 278.4 ;
         LAYER MET3 ;
         RECT  0.0 364.32 682.28 364.88 ;
         LAYER MET4 ;
         RECT  680.8 0.0 681.36 578.32 ;
         LAYER MET3 ;
         RECT  0.0 511.52 682.28 512.08 ;
         LAYER MET3 ;
         RECT  678.96 502.32 682.28 502.88 ;
         LAYER MET4 ;
         RECT  79.12 0.0 79.68 578.32 ;
         LAYER MET3 ;
         RECT  678.96 544.64 682.28 545.2 ;
         LAYER MET3 ;
         RECT  0.0 380.88 182.72 381.44 ;
         LAYER MET4 ;
         RECT  294.4 11.96 294.96 578.32 ;
         LAYER MET3 ;
         RECT  648.6 51.52 682.28 52.08 ;
         LAYER MET3 ;
         RECT  125.12 156.4 682.28 156.96 ;
         LAYER MET3 ;
         RECT  675.28 93.84 682.28 94.4 ;
         LAYER MET3 ;
         RECT  85.56 244.72 682.28 245.28 ;
         LAYER MET4 ;
         RECT  128.8 0.0 129.36 578.32 ;
         LAYER MET4 ;
         RECT  533.6 0.0 534.16 578.32 ;
         LAYER MET3 ;
         RECT  151.8 92.0 682.28 92.56 ;
         LAYER MET3 ;
         RECT  0.0 138.0 682.28 138.56 ;
         LAYER MET4 ;
         RECT  500.48 0.0 501.04 578.32 ;
         LAYER MET4 ;
         RECT  68.08 0.0 68.64 578.32 ;
         LAYER MET3 ;
         RECT  0.0 351.44 182.72 352.0 ;
         LAYER MET3 ;
         RECT  647.68 16.56 682.28 17.12 ;
         LAYER MET3 ;
         RECT  125.12 163.76 682.28 164.32 ;
         LAYER MET4 ;
         RECT  323.84 0.0 324.4 578.32 ;
         LAYER MET4 ;
         RECT  5.52 0.0 6.08 578.32 ;
         LAYER MET3 ;
         RECT  127.88 110.4 682.28 110.96 ;
         LAYER MET4 ;
         RECT  80.96 0.0 81.52 578.32 ;
         LAYER MET4 ;
         RECT  242.88 0.0 243.44 578.32 ;
         LAYER MET3 ;
         RECT  0.0 469.2 682.28 469.76 ;
         LAYER MET4 ;
         RECT  563.04 0.0 563.6 578.32 ;
         LAYER MET3 ;
         RECT  178.48 390.08 682.28 390.64 ;
         LAYER MET3 ;
         RECT  0.0 460.0 682.28 460.56 ;
         LAYER MET3 ;
         RECT  0.0 312.8 682.28 313.36 ;
         LAYER MET3 ;
         RECT  0.0 150.88 182.72 151.44 ;
         LAYER MET4 ;
         RECT  288.88 0.0 289.44 578.32 ;
         LAYER MET3 ;
         RECT  678.96 108.56 682.28 109.12 ;
         LAYER MET3 ;
         RECT  0.0 202.4 682.28 202.96 ;
         LAYER MET4 ;
         RECT  342.24 26.68 342.8 578.32 ;
         LAYER MET3 ;
         RECT  0.0 167.44 682.28 168.0 ;
         LAYER MET3 ;
         RECT  0.0 57.04 682.28 57.6 ;
         LAYER MET3 ;
         RECT  678.96 101.2 682.28 101.76 ;
         LAYER MET3 ;
         RECT  149.96 104.88 682.28 105.44 ;
         LAYER MET3 ;
         RECT  0.0 158.24 122.92 158.8 ;
         LAYER MET3 ;
         RECT  0.0 73.6 682.28 74.16 ;
         LAYER MET4 ;
         RECT  454.48 0.0 455.04 578.32 ;
         LAYER MET4 ;
         RECT  292.56 0.0 293.12 578.32 ;
         LAYER MET4 ;
         RECT  169.28 0.0 169.84 578.32 ;
         LAYER MET3 ;
         RECT  178.48 333.04 682.28 333.6 ;
         LAYER MET4 ;
         RECT  334.88 0.0 335.44 578.32 ;
         LAYER MET3 ;
         RECT  678.96 158.24 682.28 158.8 ;
         LAYER MET4 ;
         RECT  610.88 0.0 611.44 578.32 ;
         LAYER MET4 ;
         RECT  664.24 0.0 664.8 578.32 ;
         LAYER MET4 ;
         RECT  230.0 0.0 230.56 578.32 ;
         LAYER MET3 ;
         RECT  0.0 77.28 119.24 77.84 ;
         LAYER MET3 ;
         RECT  178.48 290.72 682.28 291.28 ;
         LAYER MET4 ;
         RECT  126.96 0.0 127.52 578.32 ;
         LAYER MET4 ;
         RECT  395.6 0.0 396.16 578.32 ;
         LAYER MET3 ;
         RECT  0.0 518.88 682.28 519.44 ;
         LAYER MET3 ;
         RECT  0.0 69.92 682.28 70.48 ;
         LAYER MET4 ;
         RECT  528.08 0.0 528.64 578.32 ;
         LAYER MET3 ;
         RECT  179.4 66.24 682.28 66.8 ;
         LAYER MET4 ;
         RECT  509.68 0.0 510.24 578.32 ;
         LAYER MET4 ;
         RECT  283.36 0.0 283.92 578.32 ;
         LAYER MET4 ;
         RECT  645.84 0.0 646.4 16.2 ;
         LAYER MET3 ;
         RECT  0.0 441.6 682.28 442.16 ;
         LAYER MET3 ;
         RECT  0.0 79.12 7.0 79.68 ;
         LAYER MET4 ;
         RECT  99.36 0.0 99.92 578.32 ;
         LAYER MET4 ;
         RECT  185.84 0.0 186.4 578.32 ;
         LAYER MET3 ;
         RECT  0.0 204.24 106.36 204.8 ;
         LAYER MET4 ;
         RECT  220.8 0.0 221.36 10.68 ;
         LAYER MET3 ;
         RECT  0.0 371.68 682.28 372.24 ;
         LAYER MET4 ;
         RECT  257.6 0.0 258.16 578.32 ;
         LAYER MET3 ;
         RECT  0.0 176.64 106.36 177.2 ;
         LAYER MET3 ;
         RECT  0.0 51.52 190.08 52.08 ;
         LAYER MET3 ;
         RECT  0.0 574.08 182.72 574.64 ;
         LAYER MET4 ;
         RECT  114.08 0.0 114.64 578.32 ;
         LAYER MET4 ;
         RECT  678.96 0.0 679.52 578.32 ;
         LAYER MET4 ;
         RECT  616.4 0.0 616.96 10.68 ;
         LAYER MET4 ;
         RECT  583.28 45.08 583.84 578.32 ;
         LAYER MET3 ;
         RECT  0.0 430.56 182.72 431.12 ;
         LAYER MET3 ;
         RECT  0.0 16.56 342.8 17.12 ;
         LAYER MET3 ;
         RECT  420.44 9.2 682.28 9.76 ;
         LAYER MET3 ;
         RECT  0.0 384.56 682.28 385.12 ;
         LAYER MET3 ;
         RECT  0.0 447.12 682.28 447.68 ;
         LAYER MET4 ;
         RECT  673.44 0.0 674.0 578.32 ;
         LAYER MET4 ;
         RECT  314.64 0.0 315.2 578.32 ;
         LAYER MET4 ;
         RECT  415.84 6.44 416.4 578.32 ;
         LAYER MET4 ;
         RECT  458.16 0.0 458.72 578.32 ;
         LAYER MET3 ;
         RECT  0.0 425.04 682.28 425.6 ;
         LAYER MET4 ;
         RECT  461.84 45.08 462.4 578.32 ;
         LAYER MET3 ;
         RECT  678.96 487.6 682.28 488.16 ;
         LAYER MET3 ;
         RECT  0.0 522.56 682.28 523.12 ;
         LAYER MET4 ;
         RECT  316.48 6.44 317.04 578.32 ;
         LAYER MET4 ;
         RECT  355.12 0.0 355.68 578.32 ;
         LAYER MET3 ;
         RECT  0.0 185.84 182.72 186.4 ;
         LAYER MET3 ;
         RECT  678.96 458.16 682.28 458.72 ;
         LAYER MET4 ;
         RECT  644.0 0.0 644.56 578.32 ;
         LAYER MET3 ;
         RECT  0.0 377.2 147.76 377.76 ;
         LAYER MET4 ;
         RECT  82.8 0.0 83.36 578.32 ;
         LAYER MET4 ;
         RECT  108.56 0.0 109.12 578.32 ;
         LAYER MET3 ;
         RECT  0.0 274.16 682.28 274.72 ;
         LAYER MET3 ;
         RECT  178.48 434.24 682.28 434.8 ;
         LAYER MET4 ;
         RECT  616.4 26.68 616.96 578.32 ;
         LAYER MET3 ;
         RECT  178.48 318.32 682.28 318.88 ;
         LAYER MET3 ;
         RECT  178.48 347.76 682.28 348.32 ;
         LAYER MET4 ;
         RECT  299.92 6.44 300.48 578.32 ;
         LAYER MET3 ;
         RECT  0.0 1.84 682.28 2.4 ;
         LAYER MET3 ;
         RECT  102.12 255.76 682.28 256.32 ;
         LAYER MET4 ;
         RECT  476.56 0.0 477.12 578.32 ;
         LAYER MET3 ;
         RECT  0.0 561.2 682.28 561.76 ;
         LAYER MET3 ;
         RECT  0.0 544.64 182.72 545.2 ;
         LAYER MET3 ;
         RECT  678.96 272.32 682.28 272.88 ;
         LAYER MET3 ;
         RECT  0.0 252.08 682.28 252.64 ;
         LAYER MET4 ;
         RECT  638.48 0.0 639.04 578.32 ;
         LAYER MET3 ;
         RECT  678.96 393.76 682.28 394.32 ;
         LAYER MET3 ;
         RECT  0.0 184.0 682.28 184.56 ;
         LAYER MET3 ;
         RECT  0.0 128.8 7.0 129.36 ;
         LAYER MET3 ;
         RECT  0.0 564.88 682.28 565.44 ;
         LAYER MET3 ;
         RECT  0.0 557.52 682.28 558.08 ;
         LAYER MET4 ;
         RECT  360.64 13.8 361.2 578.32 ;
         LAYER MET4 ;
         RECT  244.72 0.0 245.28 5.16 ;
         LAYER MET3 ;
         RECT  125.12 206.08 682.28 206.64 ;
         LAYER MET3 ;
         RECT  0.0 494.96 182.72 495.52 ;
         LAYER MET4 ;
         RECT  579.6 0.0 580.16 578.32 ;
         LAYER MET3 ;
         RECT  0.0 132.48 106.36 133.04 ;
         LAYER MET3 ;
         RECT  0.0 342.24 682.28 342.8 ;
         LAYER MET4 ;
         RECT  285.2 0.0 285.76 578.32 ;
         LAYER MET3 ;
         RECT  678.96 351.44 682.28 352.0 ;
         LAYER MET4 ;
         RECT  507.84 0.0 508.4 578.32 ;
         LAYER MET3 ;
         RECT  0.0 301.76 182.72 302.32 ;
         LAYER MET3 ;
         RECT  0.0 368.0 682.28 368.56 ;
         LAYER MET4 ;
         RECT  121.44 0.0 122.0 578.32 ;
         LAYER MET4 ;
         RECT  434.24 0.0 434.8 14.36 ;
         LAYER MET4 ;
         RECT  195.04 0.0 195.6 5.16 ;
         LAYER MET4 ;
         RECT  69.92 0.0 70.48 578.32 ;
         LAYER MET4 ;
         RECT  653.2 0.0 653.76 578.32 ;
         LAYER MET4 ;
         RECT  27.6 0.0 28.16 578.32 ;
         LAYER MET3 ;
         RECT  0.0 533.6 147.76 534.16 ;
         LAYER MET4 ;
         RECT  493.12 45.08 493.68 578.32 ;
         LAYER MET4 ;
         RECT  261.28 13.8 261.84 578.32 ;
         LAYER MET3 ;
         RECT  0.0 487.6 182.72 488.16 ;
         LAYER MET4 ;
         RECT  603.52 0.0 604.08 578.32 ;
         LAYER MET3 ;
         RECT  0.0 231.84 682.28 232.4 ;
         LAYER MET3 ;
         RECT  0.0 310.96 682.28 311.52 ;
         LAYER MET3 ;
         RECT  0.0 419.52 147.76 420.08 ;
         LAYER MET4 ;
         RECT  14.72 0.0 15.28 578.32 ;
         LAYER MET4 ;
         RECT  88.32 0.0 88.88 578.32 ;
         LAYER MET4 ;
         RECT  550.16 0.0 550.72 578.32 ;
         LAYER MET3 ;
         RECT  103.04 263.12 682.28 263.68 ;
         LAYER MET3 ;
         RECT  0.0 485.76 682.28 486.32 ;
         LAYER MET4 ;
         RECT  40.48 0.0 41.04 578.32 ;
         LAYER MET4 ;
         RECT  202.4 0.0 202.96 578.32 ;
         LAYER MET3 ;
         RECT  678.96 529.92 682.28 530.48 ;
         LAYER MET3 ;
         RECT  125.12 220.8 682.28 221.36 ;
         LAYER MET3 ;
         RECT  0.0 428.72 682.28 429.28 ;
         LAYER MET3 ;
         RECT  678.96 193.2 682.28 193.76 ;
         LAYER MET4 ;
         RECT  25.76 0.0 26.32 578.32 ;
         LAYER MET3 ;
         RECT  39.56 33.12 682.28 33.68 ;
         LAYER MET3 ;
         RECT  0.0 305.44 147.76 306.0 ;
         LAYER MET3 ;
         RECT  678.96 279.68 682.28 280.24 ;
         LAYER MET4 ;
         RECT  38.64 33.12 39.2 578.32 ;
         LAYER MET4 ;
         RECT  373.52 0.0 374.08 12.52 ;
         LAYER MET4 ;
         RECT  482.08 0.0 482.64 578.32 ;
         LAYER MET3 ;
         RECT  678.96 380.88 682.28 381.44 ;
         LAYER MET3 ;
         RECT  96.6 36.8 682.28 37.36 ;
         LAYER MET3 ;
         RECT  0.0 86.48 682.28 87.04 ;
         LAYER MET3 ;
         RECT  678.96 294.4 682.28 294.96 ;
         LAYER MET3 ;
         RECT  0.0 414.0 682.28 414.56 ;
         LAYER MET4 ;
         RECT  312.8 26.68 313.36 578.32 ;
         LAYER MET4 ;
         RECT  310.96 0.0 311.52 5.16 ;
         LAYER MET4 ;
         RECT  145.36 0.0 145.92 578.32 ;
         LAYER MET3 ;
         RECT  132.48 77.28 682.28 77.84 ;
         LAYER MET3 ;
         RECT  0.0 174.8 106.36 175.36 ;
         LAYER MET3 ;
         RECT  678.96 423.2 682.28 423.76 ;
         LAYER MET4 ;
         RECT  596.16 0.0 596.72 578.32 ;
         LAYER MET3 ;
         RECT  0.0 336.72 182.72 337.28 ;
         LAYER MET3 ;
         RECT  0.0 531.76 682.28 532.32 ;
         LAYER MET3 ;
         RECT  556.6 12.88 682.28 13.44 ;
         LAYER MET4 ;
         RECT  103.04 0.0 103.6 578.32 ;
         LAYER MET4 ;
         RECT  373.52 26.68 374.08 578.32 ;
         LAYER MET3 ;
         RECT  0.0 33.12 5.16 33.68 ;
         LAYER MET3 ;
         RECT  0.0 266.8 86.12 267.36 ;
         LAYER MET3 ;
         RECT  0.0 281.52 682.28 282.08 ;
         LAYER MET3 ;
         RECT  678.96 287.04 682.28 287.6 ;
         LAYER MET4 ;
         RECT  494.96 26.68 495.52 578.32 ;
         LAYER MET4 ;
         RECT  66.24 0.0 66.8 578.32 ;
         LAYER MET3 ;
         RECT  0.0 520.72 147.76 521.28 ;
         LAYER MET3 ;
         RECT  16.56 62.56 682.28 63.12 ;
         LAYER MET3 ;
         RECT  0.0 491.28 147.76 491.84 ;
         LAYER MET3 ;
         RECT  0.0 482.08 682.28 482.64 ;
         LAYER MET4 ;
         RECT  53.36 0.0 53.92 578.32 ;
         LAYER MET4 ;
         RECT  452.64 0.0 453.2 578.32 ;
         LAYER MET4 ;
         RECT  189.52 45.08 190.08 578.32 ;
         LAYER MET4 ;
         RECT  594.32 0.0 594.88 578.32 ;
         LAYER MET3 ;
         RECT  0.0 493.12 682.28 493.68 ;
         LAYER MET4 ;
         RECT  1.84 135.24 2.4 578.32 ;
         LAYER MET4 ;
         RECT  220.8 26.68 221.36 578.32 ;
         LAYER MET4 ;
         RECT  77.28 0.0 77.84 578.32 ;
         LAYER MET3 ;
         RECT  678.96 366.16 682.28 366.72 ;
         LAYER MET4 ;
         RECT  23.92 0.0 24.48 578.32 ;
         LAYER MET3 ;
         RECT  647.68 18.4 682.28 18.96 ;
         LAYER MET3 ;
         RECT  678.96 329.36 682.28 329.92 ;
         LAYER MET4 ;
         RECT  351.44 0.0 352.0 578.32 ;
         LAYER MET3 ;
         RECT  678.96 336.72 682.28 337.28 ;
         LAYER MET3 ;
         RECT  0.0 198.72 122.92 199.28 ;
         LAYER MET4 ;
         RECT  277.84 0.0 278.4 5.16 ;
         LAYER MET4 ;
         RECT  531.76 0.0 532.32 578.32 ;
         LAYER MET4 ;
         RECT  423.2 0.0 423.76 578.32 ;
         LAYER MET4 ;
         RECT  513.36 0.0 513.92 578.32 ;
         LAYER MET3 ;
         RECT  0.0 38.64 29.08 39.2 ;
         LAYER MET3 ;
         RECT  0.0 402.96 682.28 403.52 ;
         LAYER MET4 ;
         RECT  522.56 45.08 523.12 578.32 ;
         LAYER MET3 ;
         RECT  0.0 215.28 122.92 215.84 ;
         LAYER MET4 ;
         RECT  193.2 0.0 193.76 578.32 ;
         LAYER MET4 ;
         RECT  570.4 0.0 570.96 578.32 ;
         LAYER MET4 ;
         RECT  178.48 11.96 179.04 578.32 ;
         LAYER MET3 ;
         RECT  96.6 71.76 682.28 72.32 ;
         LAYER MET4 ;
         RECT  667.92 0.0 668.48 578.32 ;
         LAYER MET3 ;
         RECT  0.0 112.24 7.0 112.8 ;
         LAYER MET3 ;
         RECT  0.0 528.08 682.28 528.64 ;
         LAYER MET4 ;
         RECT  156.4 0.0 156.96 578.32 ;
         LAYER MET3 ;
         RECT  0.0 90.16 682.28 90.72 ;
         LAYER MET3 ;
         RECT  19.32 82.8 682.28 83.36 ;
         LAYER MET4 ;
         RECT  426.88 0.0 427.44 5.16 ;
         LAYER MET4 ;
         RECT  171.12 0.0 171.68 578.32 ;
         LAYER MET4 ;
         RECT  209.76 0.0 210.32 578.32 ;
         LAYER MET4 ;
         RECT  540.96 0.0 541.52 578.32 ;
         LAYER MET3 ;
         RECT  0.0 421.36 682.28 421.92 ;
         LAYER MET3 ;
         RECT  0.0 172.96 682.28 173.52 ;
         LAYER MET3 ;
         RECT  0.0 288.88 682.28 289.44 ;
         LAYER MET4 ;
         RECT  386.4 0.0 386.96 578.32 ;
         LAYER MET4 ;
         RECT  404.8 0.0 405.36 578.32 ;
         LAYER MET3 ;
         RECT  125.12 112.24 682.28 112.8 ;
         LAYER MET3 ;
         RECT  678.96 185.84 682.28 186.4 ;
         LAYER MET4 ;
         RECT  520.72 0.0 521.28 578.32 ;
         LAYER MET4 ;
         RECT  377.2 0.0 377.76 5.16 ;
         LAYER MET3 ;
         RECT  0.0 23.92 682.28 24.48 ;
         LAYER MET3 ;
         RECT  0.0 555.68 682.28 556.24 ;
         LAYER MET3 ;
         RECT  678.96 358.8 682.28 359.36 ;
         LAYER MET4 ;
         RECT  255.76 0.0 256.32 578.32 ;
         LAYER MET3 ;
         RECT  0.0 211.6 122.92 212.16 ;
         LAYER MET4 ;
         RECT  18.4 0.0 18.96 578.32 ;
         LAYER MET3 ;
         RECT  178.48 147.2 682.28 147.76 ;
         LAYER MET3 ;
         RECT  0.0 575.92 682.28 576.48 ;
         LAYER MET3 ;
         RECT  0.0 259.44 682.28 260.0 ;
         LAYER MET3 ;
         RECT  0.0 529.92 182.72 530.48 ;
         LAYER MET4 ;
         RECT  601.68 0.0 602.24 578.32 ;
         LAYER MET3 ;
         RECT  0.0 248.4 682.28 248.96 ;
         LAYER MET3 ;
         RECT  0.0 20.24 682.28 20.8 ;
         LAYER MET4 ;
         RECT  623.76 0.0 624.32 578.32 ;
         LAYER MET3 ;
         RECT  0.0 410.32 682.28 410.88 ;
         LAYER MET4 ;
         RECT  20.24 0.0 20.8 578.32 ;
         LAYER MET4 ;
         RECT  86.48 0.0 87.04 578.32 ;
         LAYER MET3 ;
         RECT  0.0 180.32 122.92 180.88 ;
         LAYER MET4 ;
         RECT  115.92 0.0 116.48 578.32 ;
         LAYER MET3 ;
         RECT  0.0 141.68 682.28 142.24 ;
         LAYER MET3 ;
         RECT  0.0 285.2 682.28 285.76 ;
         LAYER MET4 ;
         RECT  450.8 0.0 451.36 578.32 ;
         LAYER MET3 ;
         RECT  0.0 25.76 190.08 26.32 ;
         LAYER MET3 ;
         RECT  0.0 395.6 682.28 396.16 ;
         LAYER MET3 ;
         RECT  178.48 174.8 682.28 175.36 ;
         LAYER MET3 ;
         RECT  678.96 128.8 682.28 129.36 ;
         LAYER MET3 ;
         RECT  0.0 58.88 95.32 59.44 ;
         LAYER MET4 ;
         RECT  447.12 0.0 447.68 578.32 ;
         LAYER MET3 ;
         RECT  0.0 489.44 682.28 490.0 ;
         LAYER MET3 ;
         RECT  0.0 375.36 682.28 375.92 ;
         LAYER MET3 ;
         RECT  178.48 419.52 682.28 420.08 ;
         LAYER MET3 ;
         RECT  0.0 524.4 182.72 524.96 ;
         LAYER MET3 ;
         RECT  678.96 264.96 682.28 265.52 ;
         LAYER MET3 ;
         RECT  0.0 552.0 182.72 552.56 ;
         LAYER MET3 ;
         RECT  178.48 261.28 682.28 261.84 ;
         LAYER MET3 ;
         RECT  0.0 344.08 182.72 344.64 ;
         LAYER MET3 ;
         RECT  678.96 171.12 682.28 171.68 ;
         LAYER MET3 ;
         RECT  678.96 230.0 682.28 230.56 ;
         LAYER MET3 ;
         RECT  678.96 136.16 682.28 136.72 ;
         LAYER MET3 ;
         RECT  0.0 355.12 682.28 355.68 ;
         LAYER MET3 ;
         RECT  0.0 171.12 122.92 171.68 ;
         LAYER MET3 ;
         RECT  0.0 553.84 682.28 554.4 ;
         LAYER MET3 ;
         RECT  0.0 47.84 682.28 48.4 ;
         LAYER MET3 ;
         RECT  46.92 49.68 682.28 50.24 ;
         LAYER MET3 ;
         RECT  0.0 360.64 682.28 361.2 ;
         LAYER MET3 ;
         RECT  0.0 423.2 182.72 423.76 ;
         LAYER MET4 ;
         RECT  636.64 0.0 637.2 578.32 ;
         LAYER MET3 ;
         RECT  0.0 114.08 122.92 114.64 ;
         LAYER MET3 ;
         RECT  0.0 515.2 682.28 515.76 ;
         LAYER MET3 ;
         RECT  125.12 178.48 682.28 179.04 ;
         LAYER MET4 ;
         RECT  642.16 0.0 642.72 578.32 ;
         LAYER MET4 ;
         RECT  294.4 0.0 294.96 5.16 ;
         LAYER MET3 ;
         RECT  0.0 178.48 122.92 179.04 ;
         LAYER MET4 ;
         RECT  463.68 26.68 464.24 578.32 ;
         LAYER MET3 ;
         RECT  0.0 93.84 186.4 94.4 ;
         LAYER MET3 ;
         RECT  0.0 401.12 182.72 401.68 ;
         LAYER MET3 ;
         RECT  0.0 29.44 32.76 30.0 ;
         LAYER MET3 ;
         RECT  678.96 301.76 682.28 302.32 ;
         LAYER MET3 ;
         RECT  177.56 75.44 682.28 76.0 ;
         LAYER MET4 ;
         RECT  217.12 6.44 217.68 578.32 ;
         LAYER MET3 ;
         RECT  132.48 60.72 682.28 61.28 ;
         LAYER MET3 ;
         RECT  0.0 500.48 682.28 501.04 ;
         LAYER MET4 ;
         RECT  303.6 0.0 304.16 578.32 ;
         LAYER MET3 ;
         RECT  0.0 241.04 682.28 241.6 ;
         LAYER MET3 ;
         RECT  678.96 386.4 682.28 386.96 ;
         LAYER MET4 ;
         RECT  621.92 0.0 622.48 578.32 ;
         LAYER MET3 ;
         RECT  0.0 250.24 86.12 250.8 ;
         LAYER MET4 ;
         RECT  358.8 0.0 359.36 578.32 ;
         LAYER MET3 ;
         RECT  137.08 211.6 682.28 212.16 ;
         LAYER MET3 ;
         RECT  0.0 535.44 682.28 536.0 ;
         LAYER MET3 ;
         RECT  0.0 226.32 682.28 226.88 ;
         LAYER MET4 ;
         RECT  318.32 0.0 318.88 578.32 ;
         LAYER MET3 ;
         RECT  646.76 42.32 682.28 42.88 ;
         LAYER MET4 ;
         RECT  279.68 45.08 280.24 578.32 ;
         LAYER MET4 ;
         RECT  320.16 0.0 320.72 578.32 ;
         LAYER MET4 ;
         RECT  410.32 0.0 410.88 5.16 ;
         LAYER MET3 ;
         RECT  178.48 117.76 682.28 118.32 ;
         LAYER MET3 ;
         RECT  0.0 458.16 182.72 458.72 ;
         LAYER MET4 ;
         RECT  557.52 0.0 558.08 578.32 ;
         LAYER MET3 ;
         RECT  0.0 126.96 122.92 127.52 ;
         LAYER MET4 ;
         RECT  526.24 0.0 526.8 578.32 ;
         LAYER MET4 ;
         RECT  390.08 0.0 390.64 578.32 ;
         LAYER MET4 ;
         RECT  498.64 0.0 499.2 578.32 ;
         LAYER MET4 ;
         RECT  677.12 0.0 677.68 578.32 ;
         LAYER MET4 ;
         RECT  305.44 0.0 306.0 578.32 ;
         LAYER MET3 ;
         RECT  0.0 191.36 682.28 191.92 ;
         LAYER MET3 ;
         RECT  0.0 513.36 682.28 513.92 ;
         LAYER MET3 ;
         RECT  0.0 276.0 147.76 276.56 ;
         LAYER MET4 ;
         RECT  296.24 0.0 296.8 578.32 ;
         LAYER MET4 ;
         RECT  322.0 0.0 322.56 578.32 ;
         LAYER MET4 ;
         RECT  402.96 45.08 403.52 578.32 ;
         LAYER MET3 ;
         RECT  0.0 563.04 147.76 563.6 ;
         LAYER MET3 ;
         RECT  0.0 502.32 182.72 502.88 ;
         LAYER MET3 ;
         RECT  0.0 40.48 5.16 41.04 ;
         LAYER MET3 ;
         RECT  0.0 559.36 182.72 559.92 ;
         LAYER MET4 ;
         RECT  64.4 0.0 64.96 578.32 ;
         LAYER MET4 ;
         RECT  609.04 0.0 609.6 578.32 ;
         LAYER MET3 ;
         RECT  0.0 366.16 182.72 366.72 ;
         LAYER MET3 ;
         RECT  0.0 327.52 682.28 328.08 ;
         LAYER MET3 ;
         RECT  678.96 309.12 682.28 309.68 ;
         LAYER MET3 ;
         RECT  0.0 436.08 682.28 436.64 ;
         LAYER MET3 ;
         RECT  0.0 222.64 122.92 223.2 ;
         LAYER MET4 ;
         RECT  325.68 0.0 326.24 578.32 ;
         LAYER MET3 ;
         RECT  0.0 12.88 210.32 13.44 ;
         LAYER MET4 ;
         RECT  605.36 0.0 605.92 578.32 ;
         LAYER MET4 ;
         RECT  259.44 0.0 260.0 578.32 ;
         LAYER MET4 ;
         RECT  379.04 0.0 379.6 578.32 ;
         LAYER MET3 ;
         RECT  85.56 270.48 682.28 271.04 ;
         LAYER MET3 ;
         RECT  178.48 476.56 682.28 477.12 ;
         LAYER MET4 ;
         RECT  658.72 0.0 659.28 578.32 ;
         LAYER MET3 ;
         RECT  178.48 448.96 682.28 449.52 ;
         LAYER MET4 ;
         RECT  200.56 6.44 201.12 578.32 ;
         LAYER MET3 ;
         RECT  178.48 276.0 682.28 276.56 ;
         LAYER MET4 ;
         RECT  298.08 6.44 298.64 578.32 ;
         LAYER MET4 ;
         RECT  139.84 0.0 140.4 578.32 ;
         LAYER MET4 ;
         RECT  393.76 17.48 394.32 578.32 ;
         LAYER MET3 ;
         RECT  0.0 334.88 682.28 335.44 ;
         LAYER MET3 ;
         RECT  0.0 550.16 682.28 550.72 ;
         LAYER MET4 ;
         RECT  504.16 0.0 504.72 578.32 ;
         LAYER MET4 ;
         RECT  656.88 0.0 657.44 578.32 ;
         LAYER MET4 ;
         RECT  662.4 0.0 662.96 578.32 ;
         LAYER MET4 ;
         RECT  555.68 26.68 556.24 578.32 ;
         LAYER MET4 ;
         RECT  228.16 11.96 228.72 578.32 ;
         LAYER MET4 ;
         RECT  539.12 0.0 539.68 578.32 ;
         LAYER MET3 ;
         RECT  0.0 106.72 147.76 107.28 ;
         LAYER MET4 ;
         RECT  246.56 0.0 247.12 578.32 ;
         LAYER MET3 ;
         RECT  678.96 445.28 682.28 445.84 ;
         LAYER MET4 ;
         RECT  158.24 0.0 158.8 578.32 ;
         LAYER MET3 ;
         RECT  0.0 161.92 106.36 162.48 ;
         LAYER MET3 ;
         RECT  0.0 412.16 682.28 412.72 ;
         LAYER MET3 ;
         RECT  125.12 119.6 682.28 120.16 ;
         LAYER MET4 ;
         RECT  371.68 45.08 372.24 578.32 ;
         LAYER MET3 ;
         RECT  678.96 143.52 682.28 144.08 ;
         LAYER MET4 ;
         RECT  93.84 0.0 94.4 578.32 ;
         LAYER MET4 ;
         RECT  465.52 0.0 466.08 578.32 ;
         LAYER MET4 ;
         RECT  237.36 0.0 237.92 578.32 ;
         LAYER MET3 ;
         RECT  0.0 88.32 93.48 88.88 ;
         LAYER MET4 ;
         RECT  517.04 0.0 517.6 578.32 ;
         LAYER MET3 ;
         RECT  0.0 209.76 682.28 210.32 ;
         LAYER MET3 ;
         RECT  0.0 568.56 682.28 569.12 ;
         LAYER MET4 ;
         RECT  631.12 0.0 631.68 578.32 ;
         LAYER MET3 ;
         RECT  0.0 570.4 682.28 570.96 ;
         LAYER MET3 ;
         RECT  178.48 58.88 682.28 59.44 ;
         LAYER MET3 ;
         RECT  0.0 548.32 147.76 548.88 ;
         LAYER MET3 ;
         RECT  125.12 134.32 682.28 134.88 ;
         LAYER MET3 ;
         RECT  0.0 408.48 182.72 409.04 ;
         LAYER MET4 ;
         RECT  49.68 0.0 50.24 578.32 ;
         LAYER MET4 ;
         RECT  443.44 0.0 444.0 578.32 ;
         LAYER MET4 ;
         RECT  263.12 0.0 263.68 578.32 ;
         LAYER MET4 ;
         RECT  347.76 6.44 348.32 578.32 ;
         LAYER MET4 ;
         RECT  143.52 0.0 144.08 578.32 ;
         LAYER MET4 ;
         RECT  537.28 0.0 537.84 578.32 ;
         LAYER MET3 ;
         RECT  0.0 461.84 147.76 462.4 ;
         LAYER MET3 ;
         RECT  617.32 11.04 682.28 11.6 ;
         LAYER MET3 ;
         RECT  0.0 68.08 682.28 68.64 ;
         LAYER MET3 ;
         RECT  678.96 373.52 682.28 374.08 ;
         LAYER MET3 ;
         RECT  0.0 147.2 147.76 147.76 ;
         LAYER MET4 ;
         RECT  620.08 0.0 620.64 578.32 ;
         LAYER MET3 ;
         RECT  0.0 318.32 147.76 318.88 ;
         LAYER MET4 ;
         RECT  172.96 0.0 173.52 578.32 ;
         LAYER MET4 ;
         RECT  191.36 0.0 191.92 10.68 ;
         LAYER MET4 ;
         RECT  327.52 13.8 328.08 578.32 ;
         LAYER MET4 ;
         RECT  333.04 6.44 333.6 578.32 ;
         LAYER MET3 ;
         RECT  0.0 478.4 682.28 478.96 ;
         LAYER MET4 ;
         RECT  366.16 6.44 366.72 578.32 ;
         LAYER MET3 ;
         RECT  0.0 143.52 182.72 144.08 ;
         LAYER MET3 ;
         RECT  0.0 189.52 147.76 190.08 ;
         LAYER MET3 ;
         RECT  678.96 215.28 682.28 215.84 ;
         LAYER MET4 ;
         RECT  274.16 0.0 274.72 578.32 ;
         LAYER MET4 ;
         RECT  196.88 0.0 197.44 578.32 ;
         LAYER MET4 ;
         RECT  327.52 0.0 328.08 5.16 ;
         LAYER MET3 ;
         RECT  0.0 393.76 182.72 394.32 ;
         LAYER MET4 ;
         RECT  546.48 0.0 547.04 578.32 ;
         LAYER MET4 ;
         RECT  564.88 0.0 565.44 578.32 ;
         LAYER MET3 ;
         RECT  0.0 298.08 682.28 298.64 ;
         LAYER MET3 ;
         RECT  0.0 373.52 182.72 374.08 ;
         LAYER MET4 ;
         RECT  261.28 0.0 261.84 5.16 ;
         LAYER MET3 ;
         RECT  0.0 7.36 682.28 7.92 ;
         LAYER MET3 ;
         RECT  0.0 480.24 182.72 480.8 ;
         LAYER MET3 ;
         RECT  0.0 542.8 682.28 543.36 ;
         LAYER MET3 ;
         RECT  0.0 206.08 122.92 206.64 ;
         LAYER MET4 ;
         RECT  167.44 6.44 168.0 578.32 ;
         LAYER MET4 ;
         RECT  206.08 0.0 206.64 578.32 ;
         LAYER MET4 ;
         RECT  7.36 0.0 7.92 578.32 ;
         LAYER MET3 ;
         RECT  0.0 49.68 30.0 50.24 ;
         LAYER MET4 ;
         RECT  669.76 0.0 670.32 578.32 ;
         LAYER MET3 ;
         RECT  678.96 552.0 682.28 552.56 ;
         LAYER MET4 ;
         RECT  207.92 0.0 208.48 578.32 ;
         LAYER MET3 ;
         RECT  678.96 465.52 682.28 466.08 ;
         LAYER MET4 ;
         RECT  340.4 45.08 340.96 578.32 ;
         LAYER MET4 ;
         RECT  414.0 6.44 414.56 578.32 ;
         LAYER MET3 ;
         RECT  0.0 356.96 682.28 357.52 ;
         LAYER MET3 ;
         RECT  0.0 439.76 682.28 440.32 ;
         LAYER MET4 ;
         RECT  309.12 45.08 309.68 578.32 ;
         LAYER MET3 ;
         RECT  678.96 537.28 682.28 537.84 ;
         LAYER MET3 ;
         RECT  0.0 196.88 122.92 197.44 ;
         LAYER MET4 ;
         RECT  47.84 0.0 48.4 578.32 ;
         LAYER MET4 ;
         RECT  132.48 0.0 133.04 578.32 ;
         LAYER MET3 ;
         RECT  0.0 338.56 682.28 339.12 ;
         LAYER MET3 ;
         RECT  178.48 161.92 682.28 162.48 ;
         LAYER MET3 ;
         RECT  0.0 268.64 682.28 269.2 ;
         LAYER MET3 ;
         RECT  0.0 347.76 147.76 348.32 ;
         LAYER MET4 ;
         RECT  660.56 0.0 661.12 578.32 ;
         LAYER MET3 ;
         RECT  0.0 237.36 83.36 237.92 ;
         LAYER MET3 ;
         RECT  0.0 566.72 182.72 567.28 ;
         LAYER MET3 ;
         RECT  0.0 200.56 122.92 201.12 ;
         LAYER MET3 ;
         RECT  0.0 353.28 682.28 353.84 ;
         LAYER MET3 ;
         RECT  678.96 509.68 682.28 510.24 ;
         LAYER MET3 ;
         RECT  0.0 437.92 182.72 438.48 ;
         LAYER MET3 ;
         RECT  0.0 417.68 682.28 418.24 ;
         LAYER MET3 ;
         RECT  0.0 426.88 682.28 427.44 ;
         LAYER MET4 ;
         RECT  345.92 0.0 346.48 578.32 ;
         LAYER MET3 ;
         RECT  678.96 180.32 682.28 180.88 ;
         LAYER MET4 ;
         RECT  252.08 26.68 252.64 578.32 ;
         LAYER MET4 ;
         RECT  180.32 0.0 180.88 578.32 ;
         LAYER MET3 ;
         RECT  0.0 53.36 93.48 53.92 ;
         LAYER MET4 ;
         RECT  397.44 0.0 398.0 578.32 ;
         LAYER MET4 ;
         RECT  51.52 0.0 52.08 578.32 ;
         LAYER MET4 ;
         RECT  649.52 0.0 650.08 578.32 ;
         LAYER MET3 ;
         RECT  0.0 345.92 682.28 346.48 ;
         LAYER MET3 ;
         RECT  0.0 290.72 147.76 291.28 ;
         LAYER MET4 ;
         RECT  152.72 0.0 153.28 578.32 ;
         LAYER MET4 ;
         RECT  412.16 0.0 412.72 578.32 ;
         LAYER MET3 ;
         RECT  0.0 397.44 682.28 398.0 ;
         LAYER MET3 ;
         RECT  0.0 434.24 147.76 434.8 ;
         LAYER MET4 ;
         RECT  329.36 0.0 329.92 578.32 ;
         LAYER MET3 ;
         RECT  98.44 228.16 682.28 228.72 ;
         LAYER MET4 ;
         RECT  575.92 0.0 576.48 578.32 ;
         LAYER MET4 ;
         RECT  307.28 0.0 307.84 578.32 ;
         LAYER MET4 ;
         RECT  264.96 0.0 265.52 578.32 ;
         LAYER MET4 ;
         RECT  174.8 0.0 175.36 578.32 ;
         LAYER MET4 ;
         RECT  154.56 0.0 155.12 578.32 ;
         LAYER MET3 ;
         RECT  178.48 461.84 682.28 462.4 ;
         LAYER MET4 ;
         RECT  55.2 0.0 55.76 578.32 ;
         LAYER MET4 ;
         RECT  213.44 0.0 214.0 578.32 ;
         LAYER MET3 ;
         RECT  33.12 40.48 682.28 41.04 ;
         LAYER MET4 ;
         RECT  388.24 0.0 388.8 578.32 ;
         LAYER MET3 ;
         RECT  0.0 362.48 147.76 363.04 ;
         LAYER MET3 ;
         RECT  0.0 257.6 182.72 258.16 ;
         LAYER MET4 ;
         RECT  437.92 0.0 438.48 578.32 ;
         LAYER MET3 ;
         RECT  0.0 432.4 682.28 432.96 ;
         LAYER MET3 ;
         RECT  178.48 563.04 682.28 563.6 ;
         LAYER MET4 ;
         RECT  566.72 0.0 567.28 578.32 ;
         LAYER MET4 ;
         RECT  612.72 0.0 613.28 578.32 ;
         LAYER MET3 ;
         RECT  427.8 3.68 682.28 4.24 ;
         LAYER MET3 ;
         RECT  178.48 204.24 682.28 204.8 ;
         LAYER MET3 ;
         RECT  0.0 379.04 682.28 379.6 ;
         LAYER MET3 ;
         RECT  0.0 540.96 682.28 541.52 ;
         LAYER MET4 ;
         RECT  233.68 0.0 234.24 578.32 ;
         LAYER MET4 ;
         RECT  592.48 0.0 593.04 578.32 ;
         LAYER MET4 ;
         RECT  287.04 0.0 287.6 578.32 ;
         LAYER MET4 ;
         RECT  535.44 0.0 536.0 578.32 ;
         LAYER MET4 ;
         RECT  651.36 0.0 651.92 578.32 ;
         LAYER MET3 ;
         RECT  0.0 123.28 682.28 123.84 ;
         LAYER MET4 ;
         RECT  401.12 45.08 401.68 578.32 ;
         LAYER MET4 ;
         RECT  268.64 0.0 269.2 578.32 ;
         LAYER MET3 ;
         RECT  0.0 358.8 182.72 359.36 ;
         LAYER MET3 ;
         RECT  0.0 104.88 147.76 105.44 ;
         LAYER MET4 ;
         RECT  71.76 0.0 72.32 578.32 ;
         LAYER MET3 ;
         RECT  0.0 3.68 95.32 4.24 ;
         LAYER MET3 ;
         RECT  0.0 465.52 182.72 466.08 ;
         LAYER MET4 ;
         RECT  312.8 0.0 313.36 12.52 ;
         LAYER MET4 ;
         RECT  439.76 0.0 440.32 578.32 ;
         LAYER MET4 ;
         RECT  561.2 0.0 561.76 578.32 ;
         LAYER MET4 ;
         RECT  204.24 0.0 204.8 578.32 ;
         LAYER MET3 ;
         RECT  0.0 450.8 682.28 451.36 ;
         LAYER MET3 ;
         RECT  0.0 349.6 682.28 350.16 ;
         LAYER MET3 ;
         RECT  0.0 224.48 682.28 225.04 ;
         LAYER MET3 ;
         RECT  0.0 314.64 182.72 315.2 ;
         LAYER MET3 ;
         RECT  0.0 476.56 147.76 477.12 ;
         LAYER MET3 ;
         RECT  678.96 237.36 682.28 237.92 ;
         LAYER MET3 ;
         RECT  0.0 391.92 682.28 392.48 ;
         LAYER MET3 ;
         RECT  0.0 18.4 425.6 18.96 ;
         LAYER MET3 ;
         RECT  40.48 79.12 682.28 79.68 ;
         LAYER MET4 ;
         RECT  362.48 0.0 363.04 578.32 ;
         LAYER MET3 ;
         RECT  0.0 115.92 682.28 116.48 ;
         LAYER MET4 ;
         RECT  369.84 45.08 370.4 578.32 ;
         LAYER MET4 ;
         RECT  434.24 26.68 434.8 578.32 ;
         LAYER MET4 ;
         RECT  218.96 45.08 219.52 578.32 ;
         LAYER MET3 ;
         RECT  0.0 539.12 682.28 539.68 ;
         LAYER MET4 ;
         RECT  22.08 0.0 22.64 578.32 ;
         LAYER MET3 ;
         RECT  0.0 103.04 682.28 103.6 ;
         LAYER MET4 ;
         RECT  101.2 0.0 101.76 578.32 ;
         LAYER MET3 ;
         RECT  0.0 218.96 106.36 219.52 ;
         LAYER MET3 ;
         RECT  178.48 189.52 682.28 190.08 ;
         LAYER MET4 ;
         RECT  472.88 0.0 473.44 578.32 ;
         LAYER MET3 ;
         RECT  135.24 196.88 682.28 197.44 ;
         LAYER MET3 ;
         RECT  0.0 452.64 182.72 453.2 ;
         LAYER MET3 ;
         RECT  0.0 130.64 682.28 131.2 ;
         LAYER MET4 ;
         RECT  195.04 11.96 195.6 578.32 ;
         LAYER MET4 ;
         RECT  640.32 0.0 640.88 578.32 ;
         LAYER MET3 ;
         RECT  0.0 145.36 682.28 145.92 ;
         LAYER MET3 ;
         RECT  0.0 443.44 682.28 444.0 ;
         LAYER MET4 ;
         RECT  110.4 0.0 110.96 578.32 ;
         LAYER MET4 ;
         RECT  599.84 0.0 600.4 578.32 ;
         LAYER MET3 ;
         RECT  678.96 524.4 682.28 524.96 ;
         LAYER MET4 ;
         RECT  60.72 0.0 61.28 578.32 ;
         LAYER MET3 ;
         RECT  178.48 520.72 682.28 521.28 ;
         LAYER MET4 ;
         RECT  84.64 0.0 85.2 578.32 ;
         LAYER MET4 ;
         RECT  430.56 45.08 431.12 578.32 ;
         LAYER MET4 ;
         RECT  211.6 13.8 212.16 578.32 ;
         LAYER MET4 ;
         RECT  655.04 0.0 655.6 578.32 ;
         LAYER MET3 ;
         RECT  0.0 195.04 682.28 195.6 ;
         LAYER MET3 ;
         RECT  0.0 445.28 182.72 445.84 ;
         LAYER MET4 ;
         RECT  97.52 0.0 98.08 578.32 ;
         LAYER MET4 ;
         RECT  252.08 0.0 252.64 10.68 ;
         LAYER MET4 ;
         RECT  460.0 0.0 460.56 578.32 ;
         LAYER MET4 ;
         RECT  281.52 26.68 282.08 578.32 ;
         LAYER MET3 ;
         RECT  0.0 60.72 119.24 61.28 ;
         LAYER MET4 ;
         RECT  629.28 0.0 629.84 578.32 ;
         LAYER MET3 ;
         RECT  0.0 299.92 682.28 300.48 ;
         LAYER MET3 ;
         RECT  678.96 517.04 682.28 517.6 ;
         LAYER MET3 ;
         RECT  0.0 287.04 182.72 287.6 ;
         LAYER MET4 ;
         RECT  270.48 0.0 271.04 578.32 ;
         LAYER MET4 ;
         RECT  62.56 0.0 63.12 578.32 ;
         LAYER MET3 ;
         RECT  0.0 316.48 682.28 317.04 ;
         LAYER MET3 ;
         RECT  0.0 119.6 122.92 120.16 ;
         LAYER MET3 ;
         RECT  0.0 388.24 682.28 388.8 ;
         LAYER MET3 ;
         RECT  0.0 456.32 682.28 456.88 ;
         LAYER MET4 ;
         RECT  474.72 0.0 475.28 578.32 ;
         LAYER MET3 ;
         RECT  0.0 55.2 682.28 55.76 ;
         LAYER MET3 ;
         RECT  133.4 169.28 682.28 169.84 ;
         LAYER MET3 ;
         RECT  0.0 95.68 7.0 96.24 ;
         LAYER MET4 ;
         RECT  483.92 0.0 484.48 578.32 ;
         LAYER MET4 ;
         RECT  614.56 45.08 615.12 578.32 ;
         LAYER MET4 ;
         RECT  182.16 0.0 182.72 578.32 ;
         LAYER MET3 ;
         RECT  0.0 62.56 7.0 63.12 ;
         LAYER MET4 ;
         RECT  471.04 0.0 471.6 578.32 ;
         LAYER MET3 ;
         RECT  0.0 139.84 682.28 140.4 ;
         LAYER MET4 ;
         RECT  502.32 0.0 502.88 578.32 ;
         LAYER MET4 ;
         RECT  627.44 0.0 628.0 578.32 ;
         LAYER MET3 ;
         RECT  16.56 95.68 682.28 96.24 ;
         LAYER MET4 ;
         RECT  377.2 15.64 377.76 578.32 ;
         LAYER MET4 ;
         RECT  58.88 0.0 59.44 578.32 ;
         LAYER MET3 ;
         RECT  0.0 110.4 122.92 110.96 ;
         LAYER MET3 ;
         RECT  0.0 14.72 276.56 15.28 ;
         LAYER MET3 ;
         RECT  678.96 165.6 682.28 166.16 ;
         LAYER MET4 ;
         RECT  494.96 0.0 495.52 14.36 ;
         LAYER MET3 ;
         RECT  149.96 106.72 682.28 107.28 ;
         LAYER MET3 ;
         RECT  0.0 454.48 682.28 455.04 ;
         LAYER MET4 ;
         RECT  161.92 0.0 162.48 578.32 ;
         LAYER MET4 ;
         RECT  360.64 0.0 361.2 5.16 ;
         LAYER MET4 ;
         RECT  176.64 0.0 177.2 578.32 ;
         LAYER MET3 ;
         RECT  0.0 320.16 682.28 320.72 ;
         LAYER MET3 ;
         RECT  0.0 404.8 147.76 405.36 ;
         LAYER MET4 ;
         RECT  441.6 0.0 442.16 578.32 ;
         LAYER MET3 ;
         RECT  0.0 463.68 682.28 464.24 ;
         LAYER MET3 ;
         RECT  96.6 53.36 682.28 53.92 ;
         LAYER MET3 ;
         RECT  0.0 325.68 682.28 326.24 ;
         LAYER MET3 ;
         RECT  0.0 22.08 682.28 22.64 ;
         LAYER MET3 ;
         RECT  678.96 559.36 682.28 559.92 ;
         LAYER MET3 ;
         RECT  0.0 5.52 115.56 6.08 ;
         LAYER MET4 ;
         RECT  675.28 0.0 675.84 578.32 ;
         LAYER MET4 ;
         RECT  542.8 0.0 543.36 578.32 ;
         LAYER MET4 ;
         RECT  253.92 0.0 254.48 578.32 ;
         LAYER MET4 ;
         RECT  119.6 0.0 120.16 578.32 ;
         LAYER MET3 ;
         RECT  0.0 483.92 682.28 484.48 ;
         LAYER MET4 ;
         RECT  647.68 0.0 648.24 578.32 ;
         LAYER MET3 ;
         RECT  0.0 213.44 122.92 214.0 ;
         LAYER MET3 ;
         RECT  0.0 156.4 122.92 156.96 ;
         LAYER MET4 ;
         RECT  73.6 0.0 74.16 578.32 ;
         LAYER MET4 ;
         RECT  57.04 0.0 57.6 578.32 ;
         LAYER MET3 ;
         RECT  0.0 323.84 682.28 324.4 ;
         LAYER MET4 ;
         RECT  239.2 0.0 239.76 578.32 ;
         LAYER MET4 ;
         RECT  448.96 0.0 449.52 578.32 ;
         LAYER MET3 ;
         RECT  0.0 71.76 93.48 72.32 ;
         LAYER MET3 ;
         RECT  178.48 548.32 682.28 548.88 ;
         LAYER MET4 ;
         RECT  3.68 0.0 4.24 578.32 ;
         LAYER MET4 ;
         RECT  529.92 0.0 530.48 578.32 ;
         LAYER MET4 ;
         RECT  666.08 0.0 666.64 578.32 ;
         LAYER MET3 ;
         RECT  0.0 149.04 682.28 149.6 ;
         LAYER MET3 ;
         RECT  0.0 34.96 22.64 35.52 ;
         LAYER MET4 ;
         RECT  344.08 17.48 344.64 578.32 ;
         LAYER MET4 ;
         RECT  515.2 0.0 515.76 578.32 ;
         LAYER MET4 ;
         RECT  487.6 0.0 488.16 578.32 ;
         LAYER MET3 ;
         RECT  0.0 46.0 682.28 46.56 ;
         LAYER MET3 ;
         RECT  678.96 257.6 682.28 258.16 ;
         LAYER MET4 ;
         RECT  382.72 6.44 383.28 578.32 ;
         LAYER MET4 ;
         RECT  598.0 0.0 598.56 578.32 ;
         LAYER MET4 ;
         RECT  106.72 0.0 107.28 578.32 ;
         LAYER MET4 ;
         RECT  331.2 0.0 331.76 578.32 ;
         LAYER MET3 ;
         RECT  0.0 27.6 119.24 28.16 ;
         LAYER MET4 ;
         RECT  92.0 0.0 92.56 578.32 ;
         LAYER MET3 ;
         RECT  0.0 303.6 682.28 304.16 ;
         LAYER MET4 ;
         RECT  104.88 0.0 105.44 578.32 ;
         LAYER MET3 ;
         RECT  0.0 340.4 682.28 340.96 ;
         LAYER MET3 ;
         RECT  648.6 27.6 682.28 28.16 ;
         LAYER MET3 ;
         RECT  0.0 220.8 122.92 221.36 ;
         LAYER MET3 ;
         RECT  0.0 242.88 182.72 243.44 ;
         LAYER MET3 ;
         RECT  0.0 163.76 122.92 164.32 ;
         LAYER MET3 ;
         RECT  0.0 472.88 182.72 473.44 ;
         LAYER MET4 ;
         RECT  342.24 0.0 342.8 10.68 ;
         LAYER MET3 ;
         RECT  0.0 331.2 682.28 331.76 ;
         LAYER MET3 ;
         RECT  678.96 207.92 682.28 208.48 ;
         LAYER MET4 ;
         RECT  272.32 0.0 272.88 578.32 ;
         LAYER MET4 ;
         RECT  356.96 0.0 357.52 578.32 ;
         LAYER MET3 ;
         RECT  178.48 377.2 682.28 377.76 ;
         LAYER MET4 ;
         RECT  244.72 13.8 245.28 578.32 ;
         LAYER MET4 ;
         RECT  518.88 0.0 519.44 578.32 ;
         LAYER MET4 ;
         RECT  491.28 0.0 491.84 578.32 ;
         LAYER MET3 ;
         RECT  0.0 399.28 682.28 399.84 ;
         LAYER MET4 ;
         RECT  125.12 0.0 125.68 578.32 ;
         LAYER MET4 ;
         RECT  467.36 0.0 467.92 578.32 ;
         LAYER MET4 ;
         RECT  338.56 0.0 339.12 578.32 ;
         LAYER MET4 ;
         RECT  574.08 0.0 574.64 578.32 ;
         LAYER MET4 ;
         RECT  548.32 0.0 548.88 578.32 ;
         LAYER MET3 ;
         RECT  678.96 415.84 682.28 416.4 ;
         LAYER MET3 ;
         RECT  178.48 362.48 682.28 363.04 ;
         LAYER MET4 ;
         RECT  577.76 0.0 578.32 578.32 ;
         LAYER MET3 ;
         RECT  678.96 150.88 682.28 151.44 ;
         LAYER MET3 ;
         RECT  0.0 264.96 83.36 265.52 ;
         LAYER MET3 ;
         RECT  0.0 121.44 122.92 122.0 ;
         LAYER MET4 ;
         RECT  277.84 15.64 278.4 578.32 ;
         LAYER MET4 ;
         RECT  506.0 0.0 506.56 578.32 ;
         LAYER MET4 ;
         RECT  425.04 0.0 425.6 578.32 ;
         LAYER MET3 ;
         RECT  556.6 14.72 682.28 15.28 ;
         LAYER MET3 ;
         RECT  678.96 437.92 682.28 438.48 ;
         LAYER MET3 ;
         RECT  131.56 154.56 682.28 155.12 ;
         LAYER MET3 ;
         RECT  0.0 244.72 83.36 245.28 ;
         LAYER MET3 ;
         RECT  0.0 382.72 682.28 383.28 ;
         LAYER MET4 ;
         RECT  559.36 0.0 559.92 578.32 ;
         LAYER MET4 ;
         RECT  419.52 0.0 420.08 578.32 ;
         LAYER MET3 ;
         RECT  678.96 430.56 682.28 431.12 ;
         LAYER MET3 ;
         RECT  0.0 294.4 182.72 294.96 ;
         LAYER MET4 ;
         RECT  586.96 0.0 587.52 578.32 ;
         LAYER MET3 ;
         RECT  0.0 546.48 682.28 547.04 ;
         LAYER MET4 ;
         RECT  406.64 0.0 407.2 578.32 ;
         LAYER MET4 ;
         RECT  485.76 0.0 486.32 578.32 ;
         LAYER MET4 ;
         RECT  95.68 0.0 96.24 578.32 ;
         LAYER MET3 ;
         RECT  125.12 126.96 682.28 127.52 ;
         LAYER MET4 ;
         RECT  645.84 26.68 646.4 578.32 ;
         LAYER MET3 ;
         RECT  178.48 491.28 682.28 491.84 ;
         LAYER MET4 ;
         RECT  421.36 0.0 421.92 578.32 ;
         LAYER MET3 ;
         RECT  96.6 88.32 682.28 88.88 ;
         LAYER MET3 ;
         RECT  678.96 200.56 682.28 201.12 ;
         LAYER MET3 ;
         RECT  647.68 25.76 682.28 26.32 ;
         LAYER MET4 ;
         RECT  33.12 0.0 33.68 578.32 ;
         LAYER MET4 ;
         RECT  276.0 0.0 276.56 578.32 ;
         LAYER MET4 ;
         RECT  150.88 0.0 151.44 578.32 ;
         LAYER MET4 ;
         RECT  224.48 0.0 225.04 578.32 ;
         LAYER MET4 ;
         RECT  226.32 0.0 226.88 578.32 ;
         LAYER MET3 ;
         RECT  0.0 154.56 122.92 155.12 ;
         LAYER MET4 ;
         RECT  248.4 45.08 248.96 578.32 ;
         LAYER MET4 ;
         RECT  618.24 0.0 618.8 578.32 ;
         LAYER MET4 ;
         RECT  75.44 0.0 76.0 578.32 ;
         LAYER MET4 ;
         RECT  410.32 11.96 410.88 578.32 ;
         LAYER MET3 ;
         RECT  0.0 509.68 182.72 510.24 ;
         LAYER MET3 ;
         RECT  0.0 165.6 122.92 166.16 ;
         LAYER MET4 ;
         RECT  222.64 0.0 223.2 578.32 ;
         LAYER MET4 ;
         RECT  478.4 0.0 478.96 578.32 ;
         LAYER MET4 ;
         RECT  163.76 0.0 164.32 578.32 ;
         LAYER MET4 ;
         RECT  149.04 6.44 149.6 578.32 ;
         LAYER MET3 ;
         RECT  678.96 401.12 682.28 401.68 ;
         LAYER MET3 ;
         RECT  0.0 80.96 682.28 81.52 ;
         LAYER MET3 ;
         RECT  0.0 99.36 682.28 99.92 ;
         LAYER MET4 ;
         RECT  353.28 0.0 353.84 578.32 ;
         LAYER MET4 ;
         RECT  391.92 0.0 392.48 578.32 ;
         LAYER MET3 ;
         RECT  0.0 261.28 147.76 261.84 ;
         LAYER MET4 ;
         RECT  123.28 0.0 123.84 578.32 ;
         LAYER MET3 ;
         RECT  0.0 572.24 682.28 572.8 ;
         LAYER MET3 ;
         RECT  0.0 498.64 682.28 499.2 ;
         LAYER MET4 ;
         RECT  480.24 0.0 480.8 578.32 ;
         LAYER MET3 ;
         RECT  35.88 34.96 682.28 35.52 ;
         LAYER MET4 ;
         RECT  184.0 6.44 184.56 578.32 ;
         LAYER MET3 ;
         RECT  125.12 213.44 682.28 214.0 ;
         LAYER MET3 ;
         RECT  125.12 198.72 682.28 199.28 ;
         LAYER MET4 ;
         RECT  42.32 0.0 42.88 578.32 ;
         LAYER MET4 ;
         RECT  456.32 0.0 456.88 578.32 ;
         LAYER MET3 ;
         RECT  178.48 506.0 682.28 506.56 ;
         LAYER MET3 ;
         RECT  678.96 322.0 682.28 322.56 ;
         LAYER MET3 ;
         RECT  178.48 218.96 682.28 219.52 ;
         LAYER MET4 ;
         RECT  31.28 0.0 31.84 578.32 ;
         LAYER MET4 ;
         RECT  368.0 0.0 368.56 578.32 ;
         LAYER MET4 ;
         RECT  436.08 0.0 436.64 578.32 ;
         LAYER MET3 ;
         RECT  0.0 526.24 682.28 526.8 ;
         LAYER MET3 ;
         RECT  0.0 136.16 122.92 136.72 ;
         LAYER MET3 ;
         RECT  178.48 305.44 682.28 306.0 ;
         LAYER MET3 ;
         RECT  0.0 296.24 682.28 296.8 ;
         LAYER MET3 ;
         RECT  178.48 404.8 682.28 405.36 ;
         LAYER MET3 ;
         RECT  678.96 314.64 682.28 315.2 ;
         LAYER MET4 ;
         RECT  198.72 0.0 199.28 578.32 ;
         LAYER MET4 ;
         RECT  380.88 0.0 381.44 578.32 ;
         LAYER MET3 ;
         RECT  0.0 369.84 682.28 370.4 ;
         LAYER MET4 ;
         RECT  301.76 0.0 302.32 578.32 ;
         LAYER MET4 ;
         RECT  511.52 0.0 512.08 578.32 ;
         LAYER MET3 ;
         RECT  0.0 152.72 682.28 153.28 ;
         LAYER MET4 ;
         RECT  46.0 0.0 46.56 578.32 ;
         LAYER MET3 ;
         RECT  678.96 480.24 682.28 480.8 ;
         LAYER MET4 ;
         RECT  191.36 26.68 191.92 578.32 ;
         LAYER MET3 ;
         RECT  0.0 474.72 682.28 475.28 ;
         LAYER MET4 ;
         RECT  266.8 6.44 267.36 578.32 ;
         LAYER MET4 ;
         RECT  544.64 0.0 545.2 578.32 ;
         LAYER MET3 ;
         RECT  0.0 11.04 177.2 11.6 ;
         LAYER MET4 ;
         RECT  250.24 6.44 250.8 578.32 ;
         LAYER MET4 ;
         RECT  160.08 0.0 160.64 578.32 ;
         LAYER MET4 ;
         RECT  349.6 6.44 350.16 578.32 ;
         LAYER MET3 ;
         RECT  0.0 333.04 147.76 333.6 ;
         LAYER MET4 ;
         RECT  290.72 0.0 291.28 578.32 ;
         LAYER MET4 ;
         RECT  211.6 0.0 212.16 5.16 ;
         LAYER MET3 ;
         RECT  178.48 176.64 682.28 177.2 ;
         LAYER MET3 ;
         RECT  85.56 253.92 682.28 254.48 ;
         LAYER MET4 ;
         RECT  141.68 0.0 142.24 578.32 ;
         LAYER MET4 ;
         RECT  117.76 6.44 118.32 578.32 ;
         LAYER MET4 ;
         RECT  463.68 0.0 464.24 12.52 ;
         LAYER MET3 ;
         RECT  39.56 31.28 682.28 31.84 ;
         LAYER MET3 ;
         RECT  178.48 246.56 682.28 247.12 ;
         LAYER MET4 ;
         RECT  469.2 0.0 469.76 578.32 ;
         LAYER MET4 ;
         RECT  399.28 6.44 399.84 578.32 ;
         LAYER MET3 ;
         RECT  0.0 415.84 182.72 416.4 ;
         LAYER MET3 ;
         RECT  0.0 187.68 682.28 188.24 ;
         LAYER MET4 ;
         RECT  165.6 6.44 166.16 578.32 ;
         LAYER MET4 ;
         RECT  426.88 19.32 427.44 578.32 ;
         LAYER MET4 ;
         RECT  632.96 0.0 633.52 578.32 ;
         LAYER MET3 ;
         RECT  678.96 344.08 682.28 344.64 ;
         LAYER MET3 ;
         RECT  678.96 222.64 682.28 223.2 ;
         LAYER MET3 ;
         RECT  0.0 182.16 682.28 182.72 ;
         LAYER MET3 ;
         RECT  178.48 533.6 682.28 534.16 ;
         LAYER MET4 ;
         RECT  585.12 45.08 585.68 578.32 ;
         LAYER MET3 ;
         RECT  0.0 504.16 682.28 504.72 ;
         LAYER MET4 ;
         RECT  344.08 0.0 344.64 5.16 ;
         LAYER MET4 ;
         RECT  625.6 0.0 626.16 578.32 ;
         LAYER MET4 ;
         RECT  215.28 6.44 215.84 578.32 ;
         LAYER MET4 ;
         RECT  44.16 0.0 44.72 578.32 ;
         LAYER MET3 ;
         RECT  678.96 242.88 682.28 243.44 ;
         LAYER MET4 ;
         RECT  12.88 0.0 13.44 578.32 ;
         LAYER MET3 ;
         RECT  427.8 5.52 682.28 6.08 ;
         LAYER MET3 ;
         RECT  0.0 406.64 682.28 407.2 ;
         LAYER MET3 ;
         RECT  100.28 239.2 682.28 239.76 ;
         LAYER MET4 ;
         RECT  489.44 0.0 490.0 578.32 ;
         LAYER MET4 ;
         RECT  187.68 45.08 188.24 578.32 ;
         LAYER MET4 ;
         RECT  178.48 0.0 179.04 5.16 ;
         LAYER MET4 ;
         RECT  524.4 45.08 524.96 578.32 ;
         LAYER MET4 ;
         RECT  147.2 0.0 147.76 578.32 ;
         LAYER MET4 ;
         RECT  607.2 0.0 607.76 578.32 ;
         LAYER MET4 ;
         RECT  445.28 0.0 445.84 578.32 ;
         LAYER MET3 ;
         RECT  0.0 506.0 147.76 506.56 ;
      END
   END gnd
   OBS
   LAYER  MET1 ;
      RECT  0.0 0.0 682.28 578.32 ;
   LAYER  MET2 ;
      RECT  0.0 0.0 682.28 578.32 ;
   LAYER  MET3 ;
      RECT  0.0 578.12 2.2 578.32 ;
      RECT  2.2 578.12 86.84 578.32 ;
      RECT  86.84 578.12 682.28 578.32 ;
      RECT  123.64 206.28 124.4 208.28 ;
      RECT  123.64 169.48 124.4 171.48 ;
      RECT  5.88 40.84 26.12 42.52 ;
      RECT  49.88 42.68 646.04 43.44 ;
      RECT  26.12 42.52 43.44 42.68 ;
      RECT  26.12 42.68 43.44 43.44 ;
      RECT  43.44 42.68 49.88 43.44 ;
      RECT  123.64 154.76 124.4 154.92 ;
      RECT  123.64 154.92 124.4 156.76 ;
      RECT  123.64 156.76 124.4 158.44 ;
      RECT  123.64 204.6 124.4 206.28 ;
      RECT  277.28 11.4 426.32 13.08 ;
      RECT  123.64 118.12 124.4 119.8 ;
      RECT  123.64 119.8 124.4 119.96 ;
      RECT  123.64 119.96 124.4 121.8 ;
      RECT  79.48 228.52 86.84 229.28 ;
      RECT  116.28 4.04 177.92 5.72 ;
      RECT  86.84 237.72 99.56 239.4 ;
      RECT  123.64 110.76 124.4 112.44 ;
      RECT  123.64 112.44 124.4 112.6 ;
      RECT  123.64 112.6 124.4 114.44 ;
      RECT  84.08 237.72 86.84 239.4 ;
      RECT  86.84 263.48 88.52 265.16 ;
      RECT  84.08 263.48 86.84 265.16 ;
      RECT  23.36 33.32 38.84 33.48 ;
      RECT  88.52 263.48 102.32 265.16 ;
      RECT  426.32 13.08 495.16 14.92 ;
      RECT  426.32 14.92 495.16 15.08 ;
      RECT  426.32 15.08 495.16 16.76 ;
      RECT  426.32 16.76 495.16 16.92 ;
      RECT  426.32 16.92 495.16 18.6 ;
      RECT  495.16 16.92 646.96 18.6 ;
      RECT  26.12 43.44 95.88 44.36 ;
      RECT  26.12 44.36 95.88 44.52 ;
      RECT  95.88 43.44 646.04 44.36 ;
      RECT  0.0 0.0 2.2 0.2 ;
      RECT  2.2 0.0 96.04 0.2 ;
      RECT  96.04 0.0 119.96 0.2 ;
      RECT  119.96 0.0 680.08 0.2 ;
      RECT  680.08 0.0 682.28 0.2 ;
      RECT  177.92 4.04 416.04 5.72 ;
      RECT  177.92 5.72 416.04 5.88 ;
      RECT  116.28 3.88 416.04 4.04 ;
      RECT  211.04 11.4 277.28 13.08 ;
      RECT  123.64 75.8 131.76 77.48 ;
      RECT  426.32 11.4 525.52 13.08 ;
      RECT  495.16 13.08 525.52 13.24 ;
      RECT  495.16 13.24 525.52 14.92 ;
      RECT  525.52 13.24 555.88 14.92 ;
      RECT  123.64 197.24 124.4 200.76 ;
      RECT  123.64 175.16 124.4 176.84 ;
      RECT  123.64 176.84 124.4 177.0 ;
      RECT  124.4 175.16 133.6 176.84 ;
      RECT  123.64 177.0 124.4 178.84 ;
      RECT  123.64 178.84 124.4 180.52 ;
      RECT  107.08 132.84 123.64 134.52 ;
      RECT  277.28 13.08 343.52 14.92 ;
      RECT  343.52 13.08 426.32 14.92 ;
      RECT  343.52 14.92 426.32 15.08 ;
      RECT  343.52 15.08 426.32 16.76 ;
      RECT  119.96 65.68 123.64 66.44 ;
      RECT  123.64 65.68 178.68 66.44 ;
      RECT  96.04 65.68 119.96 66.44 ;
      RECT  123.64 218.4 124.4 222.84 ;
      RECT  124.4 218.4 137.28 219.16 ;
      RECT  123.64 161.36 124.4 165.8 ;
      RECT  124.4 161.36 131.76 162.12 ;
      RECT  124.4 157.68 177.76 158.44 ;
      RECT  84.08 245.08 84.84 246.0 ;
      RECT  84.08 246.0 84.84 246.76 ;
      RECT  84.84 246.0 86.84 246.76 ;
      RECT  86.84 246.0 100.48 246.76 ;
      RECT  128.08 136.52 129.92 137.28 ;
      RECT  129.92 136.52 177.76 137.28 ;
      RECT  124.4 136.52 128.08 137.28 ;
      RECT  123.64 132.84 124.4 137.28 ;
      RECT  124.4 165.04 177.76 165.8 ;
      RECT  123.64 168.72 124.4 169.48 ;
      RECT  96.04 58.32 119.96 59.08 ;
      RECT  123.64 58.32 177.76 59.08 ;
      RECT  119.96 58.32 123.64 59.08 ;
      RECT  2.2 74.88 15.84 75.64 ;
      RECT  15.84 74.88 18.6 75.64 ;
      RECT  0.0 74.88 2.2 75.64 ;
      RECT  177.76 157.68 678.24 158.44 ;
      RECT  96.04 75.8 119.96 76.56 ;
      RECT  119.96 75.8 123.64 76.56 ;
      RECT  119.96 76.56 123.64 77.48 ;
      RECT  96.04 3.12 116.28 3.88 ;
      RECT  116.28 3.12 119.96 3.88 ;
      RECT  119.96 3.12 427.08 3.88 ;
      RECT  119.96 0.2 419.72 1.12 ;
      RECT  181.6 272.68 678.24 273.44 ;
      RECT  181.6 250.6 678.24 251.36 ;
      RECT  124.4 204.6 135.44 205.36 ;
      RECT  0.0 133.76 2.2 134.52 ;
      RECT  2.2 133.76 7.72 134.52 ;
      RECT  7.72 133.76 107.08 134.52 ;
      RECT  183.44 487.04 678.24 487.8 ;
      RECT  137.28 222.08 177.76 222.84 ;
      RECT  177.76 222.08 181.6 222.84 ;
      RECT  124.4 222.08 137.28 222.84 ;
      RECT  2.2 83.16 7.72 85.76 ;
      RECT  7.72 83.16 18.6 85.76 ;
      RECT  0.0 83.16 2.2 85.76 ;
      RECT  123.64 85.0 186.96 85.76 ;
      RECT  18.6 85.0 96.04 85.76 ;
      RECT  96.04 85.0 123.64 85.76 ;
      RECT  131.76 75.8 176.84 76.56 ;
      RECT  2.2 31.64 5.88 32.4 ;
      RECT  5.88 31.64 38.84 32.4 ;
      RECT  5.88 32.4 38.84 33.32 ;
      RECT  183.44 280.04 678.24 280.8 ;
      RECT  183.44 494.4 678.24 495.16 ;
      RECT  23.36 39.92 29.8 40.68 ;
      RECT  2.2 91.44 7.72 92.2 ;
      RECT  7.72 91.44 18.6 92.2 ;
      RECT  0.0 91.44 2.2 92.2 ;
      RECT  123.64 171.48 124.4 172.24 ;
      RECT  124.4 110.76 127.16 111.52 ;
      RECT  190.8 25.2 646.96 25.96 ;
      RECT  183.44 530.28 678.24 531.04 ;
      RECT  181.6 265.32 678.24 266.08 ;
      RECT  124.4 171.48 678.24 172.24 ;
      RECT  177.76 136.52 678.24 137.28 ;
      RECT  30.72 49.12 46.2 49.88 ;
      RECT  183.44 423.56 678.24 424.32 ;
      RECT  124.4 179.76 177.76 180.52 ;
      RECT  177.76 179.76 181.6 180.52 ;
      RECT  96.04 92.36 123.64 93.12 ;
      RECT  123.64 92.36 151.08 93.12 ;
      RECT  183.44 458.52 678.24 459.28 ;
      RECT  107.08 125.48 123.64 126.24 ;
      RECT  183.44 501.76 678.24 502.52 ;
      RECT  183.44 365.6 678.24 366.36 ;
      RECT  183.44 308.56 678.24 309.32 ;
      RECT  86.84 271.76 88.52 272.52 ;
      RECT  2.2 270.84 84.84 271.76 ;
      RECT  2.2 271.76 84.84 272.52 ;
      RECT  84.84 271.76 86.84 272.52 ;
      RECT  88.52 271.76 103.24 272.52 ;
      RECT  18.6 108.0 123.64 108.76 ;
      RECT  123.64 108.0 148.48 108.76 ;
      RECT  148.48 108.0 179.76 108.76 ;
      RECT  2.2 108.0 7.72 108.76 ;
      RECT  7.72 108.0 18.6 108.76 ;
      RECT  0.0 108.0 2.2 108.76 ;
      RECT  124.4 118.12 128.08 118.88 ;
      RECT  123.64 208.28 124.4 209.04 ;
      RECT  123.64 211.04 124.4 215.48 ;
      RECT  137.28 208.28 177.76 209.04 ;
      RECT  177.76 208.28 181.6 209.04 ;
      RECT  124.4 208.28 136.36 209.04 ;
      RECT  124.4 211.04 136.36 211.8 ;
      RECT  136.36 208.28 137.28 209.04 ;
      RECT  128.08 132.84 129.92 133.6 ;
      RECT  124.4 132.84 128.08 133.6 ;
      RECT  183.44 408.84 678.24 409.6 ;
      RECT  2.2 66.6 18.6 67.36 ;
      RECT  0.0 66.6 2.2 67.36 ;
      RECT  183.44 142.96 678.24 143.72 ;
      RECT  183.44 394.12 678.24 394.88 ;
      RECT  183.44 372.96 678.24 373.72 ;
      RECT  177.92 5.88 416.04 6.64 ;
      RECT  416.04 5.88 426.32 6.64 ;
      RECT  426.32 5.88 427.08 6.64 ;
      RECT  183.44 552.36 678.24 553.12 ;
      RECT  183.44 337.08 678.24 337.84 ;
      RECT  183.44 566.16 678.24 566.92 ;
      RECT  183.44 351.8 678.24 352.56 ;
      RECT  181.6 179.76 678.24 180.52 ;
      RECT  86.84 228.52 97.72 229.28 ;
      RECT  79.48 229.28 97.72 229.44 ;
      RECT  79.48 229.44 97.72 230.2 ;
      RECT  97.72 229.44 678.24 230.2 ;
      RECT  26.12 40.84 32.4 41.76 ;
      RECT  26.12 41.76 32.4 42.52 ;
      RECT  32.4 41.76 43.44 42.52 ;
      RECT  23.36 40.68 32.4 40.84 ;
      RECT  29.8 39.0 32.4 39.76 ;
      RECT  29.8 39.76 32.4 39.92 ;
      RECT  32.4 39.0 49.88 39.76 ;
      RECT  29.8 39.92 32.4 40.68 ;
      RECT  183.44 380.32 678.24 381.08 ;
      RECT  123.64 121.8 124.4 122.56 ;
      RECT  124.4 121.8 128.08 122.56 ;
      RECT  128.08 121.8 129.92 122.56 ;
      RECT  129.92 121.8 177.76 122.56 ;
      RECT  0.0 124.56 2.2 125.32 ;
      RECT  2.2 124.56 7.72 125.32 ;
      RECT  7.72 124.56 18.6 125.32 ;
      RECT  177.76 121.8 678.24 122.56 ;
      RECT  183.44 358.24 678.24 359.0 ;
      RECT  183.44 465.88 678.24 466.64 ;
      RECT  181.6 236.8 678.24 237.56 ;
      RECT  0.0 117.2 2.2 117.96 ;
      RECT  2.2 117.2 18.6 117.96 ;
      RECT  123.64 114.44 124.4 115.2 ;
      RECT  124.4 114.44 177.76 115.2 ;
      RECT  177.76 114.44 678.24 115.2 ;
      RECT  183.44 537.64 678.24 538.4 ;
      RECT  183.44 452.08 678.24 452.84 ;
      RECT  123.64 125.48 124.4 129.92 ;
      RECT  128.08 129.16 129.92 129.92 ;
      RECT  129.92 129.16 177.76 129.92 ;
      RECT  124.4 129.16 128.08 129.92 ;
      RECT  177.76 129.16 678.24 129.92 ;
      RECT  183.44 523.84 678.24 524.6 ;
      RECT  183.44 193.56 678.24 194.32 ;
      RECT  183.44 444.72 678.24 445.48 ;
      RECT  183.44 301.2 678.24 301.96 ;
      RECT  183.44 516.48 678.24 517.24 ;
      RECT  183.44 286.48 678.24 287.24 ;
      RECT  183.44 386.76 678.24 387.52 ;
      RECT  124.4 168.72 132.68 169.48 ;
      RECT  107.08 111.68 123.64 112.44 ;
      RECT  177.76 165.04 678.24 165.8 ;
      RECT  179.76 108.0 678.24 108.76 ;
      RECT  148.48 107.08 149.24 108.0 ;
      RECT  183.44 558.8 678.24 559.56 ;
      RECT  26.12 44.52 95.88 45.28 ;
      RECT  183.44 257.96 678.24 258.72 ;
      RECT  33.48 28.88 81.16 29.64 ;
      RECT  183.44 329.72 678.24 330.48 ;
      RECT  181.6 208.28 678.24 209.04 ;
      RECT  183.44 150.32 678.24 151.08 ;
      RECT  183.44 437.36 678.24 438.12 ;
      RECT  183.44 430.0 678.24 430.76 ;
      RECT  183.44 293.84 678.24 294.6 ;
      RECT  183.44 545.0 678.24 545.76 ;
      RECT  124.4 125.48 128.08 126.24 ;
      RECT  128.08 125.48 129.0 126.24 ;
      RECT  181.6 200.92 678.24 201.68 ;
      RECT  183.44 509.12 678.24 509.88 ;
      RECT  183.44 401.48 678.24 402.24 ;
      RECT  27.96 79.48 39.76 80.24 ;
      RECT  2.2 100.64 7.72 101.4 ;
      RECT  7.72 100.64 18.6 101.4 ;
      RECT  0.0 100.64 2.2 101.4 ;
      RECT  18.6 100.64 123.64 101.4 ;
      RECT  123.64 100.64 179.76 101.4 ;
      RECT  179.76 100.64 678.24 101.4 ;
      RECT  183.44 573.52 678.24 574.28 ;
      RECT  23.36 33.48 35.16 34.24 ;
      RECT  23.36 34.24 35.16 35.16 ;
      RECT  35.16 33.48 38.84 34.24 ;
      RECT  124.4 214.72 137.28 215.48 ;
      RECT  137.28 214.72 181.6 215.48 ;
      RECT  181.6 214.72 678.24 215.48 ;
      RECT  124.4 197.24 134.52 198.0 ;
      RECT  183.44 322.36 678.24 323.12 ;
      RECT  183.44 315.0 678.24 315.76 ;
      RECT  123.64 154.0 124.4 154.76 ;
      RECT  124.4 154.0 130.84 154.76 ;
      RECT  183.44 480.6 678.24 481.36 ;
      RECT  183.44 473.24 678.24 474.0 ;
      RECT  2.2 254.28 84.84 255.2 ;
      RECT  2.2 255.2 84.84 255.96 ;
      RECT  84.84 255.2 86.84 255.96 ;
      RECT  86.84 255.2 101.4 255.96 ;
      RECT  183.44 415.28 678.24 416.04 ;
      RECT  183.44 186.2 678.24 186.96 ;
      RECT  181.6 222.08 678.24 222.84 ;
      RECT  183.44 243.24 678.24 244.0 ;
   LAYER  MET4 ;
      RECT  0.0 2.2 0.2 85.0 ;
      RECT  0.0 85.0 0.2 578.32 ;
      RECT  0.0 0.0 0.2 2.2 ;
      RECT  370.2 5.88 371.88 13.24 ;
      RECT  370.2 2.2 371.88 5.88 ;
      RECT  583.64 5.88 585.32 25.96 ;
      RECT  583.64 25.96 585.32 44.36 ;
      RECT  522.92 5.88 524.6 25.96 ;
      RECT  583.64 2.2 585.32 5.88 ;
      RECT  585.32 16.92 585.48 25.96 ;
      RECT  311.16 13.24 311.32 14.92 ;
      RECT  311.32 13.24 313.0 14.92 ;
      RECT  309.48 5.88 311.16 13.24 ;
      RECT  309.48 13.24 311.16 14.92 ;
      RECT  432.6 15.08 434.44 25.96 ;
      RECT  370.2 13.24 371.88 44.36 ;
      RECT  188.04 2.2 189.72 5.88 ;
      RECT  188.04 5.88 189.72 11.4 ;
      RECT  188.04 11.4 189.72 44.36 ;
      RECT  522.92 25.96 524.6 44.36 ;
      RECT  614.92 11.4 616.6 25.96 ;
      RECT  0.2 85.0 2.04 134.52 ;
      RECT  401.48 5.88 403.16 11.4 ;
      RECT  401.48 11.4 403.16 25.96 ;
      RECT  401.48 2.2 403.16 5.72 ;
      RECT  401.48 5.72 403.16 5.88 ;
      RECT  493.32 15.08 493.48 25.96 ;
      RECT  493.48 15.08 495.16 25.96 ;
      RECT  522.92 2.2 524.6 5.88 ;
      RECT  165.96 2.2 167.64 5.72 ;
      RECT  215.64 2.2 217.32 5.72 ;
      RECT  364.68 2.2 366.36 5.72 ;
      RECT  348.12 2.2 349.8 5.72 ;
      RECT  430.92 2.2 432.6 5.72 ;
      RECT  430.92 5.72 432.6 5.88 ;
      RECT  430.92 5.88 432.6 25.96 ;
      RECT  430.92 25.96 432.6 44.36 ;
      RECT  414.36 2.2 416.04 5.72 ;
      RECT  298.44 2.2 300.12 5.72 ;
      RECT  401.48 25.96 403.16 44.36 ;
      RECT  554.2 13.24 555.88 25.96 ;
      RECT  37.16 2.2 38.84 32.4 ;
      RECT  371.88 13.24 373.72 25.96 ;
      RECT  189.88 11.4 191.56 25.96 ;
      RECT  189.72 11.4 189.88 25.96 ;
      RECT  312.24 14.92 313.0 25.96 ;
      RECT  376.64 5.88 377.4 13.24 ;
      RECT  376.64 13.24 377.4 14.92 ;
      RECT  409.76 5.88 410.52 11.24 ;
      RECT  682.08 0.0 682.28 2.2 ;
      RECT  682.08 2.2 682.28 5.88 ;
      RECT  682.08 5.88 682.28 578.32 ;
      RECT  244.16 5.88 244.92 11.4 ;
      RECT  244.16 11.4 244.92 13.08 ;
      RECT  293.84 5.88 294.6 11.24 ;
      RECT  281.88 2.2 282.64 5.88 ;
      RECT  281.88 5.88 282.64 13.24 ;
      RECT  281.88 13.24 282.64 25.96 ;
      RECT  194.48 5.88 195.24 11.24 ;
      RECT  211.04 5.88 211.8 13.08 ;
      RECT  403.16 11.4 404.08 25.96 ;
      RECT  360.08 5.88 360.84 13.08 ;
      RECT  524.6 11.4 525.52 25.96 ;
      RECT  326.96 5.88 327.72 13.08 ;
      RECT  260.72 5.88 261.48 11.4 ;
      RECT  260.72 11.4 261.48 13.08 ;
      RECT  464.04 13.24 464.8 25.96 ;
      RECT  266.24 2.2 267.0 5.72 ;
      RECT  232.2 2.2 232.96 5.72 ;
      RECT  183.44 2.2 184.2 5.72 ;
      RECT  177.92 5.88 178.68 11.24 ;
      RECT  646.2 16.92 646.96 25.96 ;
      RECT  342.6 13.24 343.36 16.76 ;
      RECT  342.6 16.76 343.36 25.96 ;
      RECT  343.36 13.24 344.28 16.76 ;
      RECT  342.6 11.4 343.52 13.24 ;
      RECT  343.52 5.88 344.28 11.4 ;
      RECT  343.52 11.4 344.28 13.24 ;
      RECT  492.56 5.88 493.32 15.08 ;
      RECT  492.56 15.08 493.32 44.36 ;
      RECT  492.56 2.2 493.32 5.88 ;
      RECT  426.32 5.88 427.08 18.6 ;
      RECT  585.48 16.92 586.24 25.96 ;
      RECT  277.28 5.88 278.04 13.24 ;
      RECT  277.28 13.24 278.04 14.92 ;
      RECT  149.4 2.2 150.16 5.72 ;
      RECT  227.6 5.88 228.36 11.24 ;
      RECT  221.16 13.24 221.92 25.96 ;
      RECT  221.16 11.4 221.92 13.24 ;
      RECT  393.2 5.88 393.96 16.76 ;
      RECT  200.0 2.2 200.76 5.72 ;
      RECT  251.52 11.4 252.28 13.24 ;
      RECT  251.52 13.24 252.28 25.96 ;
      RECT  248.76 5.88 249.52 11.4 ;
      RECT  248.76 2.2 249.52 5.72 ;
      RECT  248.76 5.72 249.52 5.88 ;
      RECT  249.52 2.2 250.44 5.72 ;
      RECT  248.76 11.4 249.52 13.08 ;
      RECT  248.76 13.08 249.52 13.24 ;
      RECT  248.76 13.24 249.52 25.96 ;
      RECT  248.76 25.96 249.52 44.36 ;
   END
END    sram_1rw0r0w_16_512_lapis20
END    LIBRARY
